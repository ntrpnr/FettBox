PK   D�LU����R  �>    cirkitFile.json�}�r%���881����~�?�{c[
�;�Iqu��"{�l��h_f�i�sx�<�BU��,���a��, �!�Hd��������f�������w�oo.>���x�����_^��������|�w�������o�{����knS�����1̊&0�ٖE7t�t�ť��������o/ϧ ��N�1`)�Dc�R�;�ƀ��w:Qx���~�������5F[�<g�1����,�f0\�Ƅf����T��7\ءgB��i#��4AI��	�$츾kt����w���7��[T�%���w��C�]`�#;�Н���K��<V�=���w��D�=�W]���H=V���!P���l��֎���D�-��x3K(L�1��c;���������y��'P��t����8�{�m/fl���>4]`�G�t+�&��r���{���(�:�@3���t�Z_�*���h_0�i!J��8�8o�F߰Fņ�֊8��1N���<�}����_ ,>��1`)�9w�K�Ϲ}@x�2�}1�\O�tpHy������'Ā��g
�j!X�,�� $����@{�[ ��I���U<���u�(�Z~�愢��y��Gb>
���U�T�
k��B�&�P��
4�d��
4���V�I$� �DB���h	^g�I��!�Q�u���l4	��c4
,	��H�(�S�ugA����������0���������R���n�?#�	Zt�]Z�hy'hyG�NТK�O�;I�;Rt��)Z�)Zޑ����N��N����E�w��w��w��-:�������#E'h��坣�):A���<-�<-�H�	Zt|hyhyG�NТ�����1�gA�O��'����.��b�B;��à�'���S�1����A!T�U�a���"m?���J9�[��B�zb�_>j"]b'�� ƗɈ�G�������5��u�uH�$gM�k��F.u3��s���A�������&1��}Z|�_>%���C�O�����#�yh�	b|�$�x[����'���3tb�{=��1�|�O�?�s�b�G�Hbׅ� Ɨo\��u��'���"��#v]h�	b|��1���Z|�_��C�?b��� Ɨo�����'���;Q�]G�[��v�ľK�7:z�m�F�W�����?{G�^}~�h]"[���qT�5�q�i�`]`Z���%������/ޑ�Q�" [�(U��T���r���ȑ3(�Xm#pc��7�Ώ/௭?�:��~�Q�Wah�5"-��t`QX����^H�'��p�k-�i��-��]�Ǐz��G���	����8k������������ȥ�x������Z�)
)
)?
)�
)�.� )�pZ����F�i�f��B��|fL˛�����$��mⴑ����G j��c���6�ŠQ�6rD�!�6�z�5___`����~-r�MD��(>����i�����2�p_�[j��Ԃ���F�5�/\R�&����}��!{]sC@M�z]sC��E�uZآ���2,x۳!_iKJ+݀�u-&)h�Q\�LP�Q�UFx#�P�imz�lc��]��8��ڦ�F�i\��*I�T�t�%��gQ�iۤ�[�T�~���H�!�eY�+ �8�cM��6:4b�6[ٰ��N*��;��`��l�BÔo�!����	
4>�6[��֑�B�7w`�qq�P]G��f�4e����>�a���ժ�(��1��Q,G�g�Y��L,|L����^߷U�OOP���
�#�9��d3^5�2�S��_,�`�o���צ@��KKb�g�k:��:��~@jڙ#;X����d�`=��d'�:lr�Š�TZ/Ԁ���@U�WI�����*����5B$׳�nҩƩ$֮0��W�ZA��pБ�v����G�5Y�����ӭ�BB�n��#g��nc����+䬫���w�(�ș�j�%�y{m��4rҪ��B!�}�xZeb�����:�iZ���݌���g�8X}�����F#�D��z]�� ?.F�UH�׸�j���<R�5R�5R�5R������?K}&��Ut(�j�隹
���h����y��<3�i�h�а���5N����j��܂Z�m��*�U&�׈��5u�5���`��ĕK���I��&�T9z�<%��zf�T�>5���]��nx���6��Oj#�b��gZU����`Ð*^&�w�1e˜k��I�u3�:�z�u�혋�k�ʔ,ٕ�^�x)��3����[׍�&i�4RJ3�T}�Y�b��0�M�fZU��{���w�;n���_������ ��]��ke�z�u*�Wi��L�fMp��VNh=��L�����&D��>MW��J�L�ַ&o\un�uP��Қ�$.1�$zi�j�j���R��H�z�MZ�x�(]/��J�bI�ž�C�:߫��A�g8�i�jd"�Y���bT�	�Q�_���q���ֽ�i9Oz!��<���-��6�_+u�iT}F��v1kF���n�dA5\[A���m��p%�/hW�v$���HI��i��nUJ@�@='%��S�"%@	�,��}t��>��S)��;IMl@��bl3I+N��\j�a�J��+��pMJ@�g�YXۈ����>��3�eN�)'����r��3���k,XۈC
Y��X����m���������<��k?#4�5���U�H�% ް��� w�Gb�5�j���z\�f����f�ju�O�f4PH0w��`e{�ɇ����'PJ�*j�|؀�ږ?�a����r���㝺"=:��Y�7F�����J@��0]���9��5��D���O1��h�FLӵMR�>@(�ʒ�b�H)��b�8	����lb���Xum�ܶ�"�	�%�BLt��Mg$Ov������i���i�f.�L+���`L����Y���i'������w���������g���yUBt�/|�� �%$���IDD�x�)4���<�hʏ!�U�"M��dBÐtl�Cd��L�$�D�8D�
�;�Chq�"�	�ҷa�!�T�P�r�����Z���atZ�Aۺ�1HLdz[��mo�JI�in�q����Lw}P�AaE\�io�׺���*"1��oqл�s되�58��`yτ�A�7�)�A*Q�6�6"I�hy�� ����
��&9�BD4i!�4�7�=!�t�E�lvA�\S�h��&�&ӐdJ���X]�$�d��� ��4w�C��Փ�Lw�.p�Z2Ldꛊ'��(�7���5�"1�)E�h�f߇V ��dj����q 2,���$��T��>h&"J|����dz���� �D��%������9�0Q���D����$��5J�_���S�g.��*6�*6����M�:�&LÁ-��M��9�	_�Y�i8�V�	V��&�J��-��M���819UB�n�Ul����y�ɩ�u�b�|7�_LN���[`�`�q^cr��|���+ߍ��S%��X�&X�n�˘�*!_��*6���?�q��6A+�A��q���F^�Fn�6~�����x^��۠-��&���-YJ�n�~m�6�n#��x`��۠�'�4(y���	�2�Ȟ�3h&l㈉m<�MЊm��s�mx��7�	Z��|~�o���6A+�A��l��m��MЊm����,l�m�Vl�6��؆���e��۠��K���F'b�m��m��6~�&h�6h�}�mx��_�	Z��|oi�n�m�Vl�6߿چ���e��۠��ȶ��6~�&h�6h�}�mx��_�	Z��2�	���8M#���&ю���7��?���^I��-����J*���O�WR�ߗ.CE�����\
XI��N����J*�[��;�T*�~WRy��;~_����nm�b��=<kǗXK��a-��s��I�Z2���b�
|-��G���$k�Tnկ%S����^��S�����Dg�F���_��*�s֒����s��d*/i֒�<4YK�F�k�9֒��ĵ
k�T�^�]ui�X�H��?E3��E)��T�u*Tb��"��5q�vzm��L����0TWL��AQ�ĕYI�.�� *n�VQY� *aɆ�I_2�adĒ�#��e`d�4�j����t)$XЈ����Ň���[BC�RH���b��v���H�\t�adh�ʣ�W�0ad�+�גY4a���##HX|���`dw�`d�o)V�~��^�{c��b�B�%�R�,
1,q	��_XҘ%���|ɾ�e_��AT�De��QY^�E�:"ᥑ�ekFF-�k��,�sЌx{2��Z>X��Ā#C#���Ϝ���h����9�c��H�5#C#��!X�8��Z24R,+� ג��b�`G�c��]ui��`�Q�֒�����^���GD�F��p蓯�))V4�Ĳ5#CcQh)�4���b�3|q-)ֆĲ�4R�i�X�H���b����~�Z2�R��Uf�Hd:oYV������	s��DE,Y������j?��<��U?��<j�yf:�1m�eMֺ޸�I�~_����Z���^�QH2Kbz�t��X���Y��� ��(uC��&&�mx��ۖ5]�����]��De�2�C�;x���q�|�-s��NQ��Y������`�m;�bb�6B�bǢWF7^Jn�2�E,�Qژ&��L�.)�{ֻ�g�mb��DeK��C�1�aZ�5�k�I�m>���+�,b��S��JCe�QԬ	.���	�CX�����mB4�3��ݨdϔj}kr���-cQY���	Mb$�M"��Fڪ�����X/U��UB�,bi��<����9�JZjImƾ�C�:߫e, *�c�I·e"$���ΰgBEkT�l'sDe�b�aH��uZ�&�L�Fۤ(��q�ʲޕm���+��7Zǂ5�ʠ�To�X�v�@T�����q *��=���ޠ��7��,tI���5B��b� �
�Ǩ�o���
�/ *�|I��}�1XZL��j%gM�'��o��<�q���,�De�/ *�|I��0]�L�k��JV�X���N?�G����AT���l5C�,�%���d0��)Mr��>)O>Hӊsn?DE,9k *�� T��!ih������u�y�B�qp���a�FSY� T$	��}@X�[XV�z�twDE-�� �_���"_@T���t��5{Q^@��@�A��/�A���߭�&���4��<_�����As����w��4��<_����/B3��_�&%_����vN�)�	�<����}��	�����⻧��KXN@���C�KDD�	/I:$�$ADD���C�KDD�	/I:$�$ADD������4*�Nkөm2�-�7����4��t� S�T�^�`"�߂L�(A�b���o�؏T��A�7h@*D�S�a�
��ą��B�<m�Ym�MZ��M�B����~�� �B�lvA�w�iH2�ME	d���E�a"S�T�@�8;&2�ME	d����a"S�t�� S�T���`"��L�SQzHXNcX��qI�ǩ(=$,��D��%���������dz���C�rLdz\��q*J	�i0��qI��k��SS=/%�:����*։���T	��։��$(2PS%��X'��p��v@M���[`�HXN"�5UB�n�u"a9	�,�T	��։��$(2PS%��X'��p��n@M���[`�HXN"�5UB�n�u"a9	���T	��։��4�6W��Ɔ�����T�rr���������*S������6��&h�������6��&h�������6.�&h�������6n�&h�������6��&h�������6��&h�������6.�&h�������6n�&h�����<Y��/��T�rr�����/��T�rr�����Hl��LNN�����e���JXNN�����e���JXNN�����e���JXNN�����e���JXNN�����e���JXNN�����e���JXNN�����e �OBtA��T�r��R�}��J��J*��+�T�$��R�E��J���J*���+�T�֮�:"ᥑ��#��dh���j-	�=hZK�F�kφ֒����㜵d�t0���^Ҭ%C#ŵ�!k��Hq��Z2D�G3�+)VD��dP4R����Oeq��	��TG	��O�f�8a9�ʢ~ ','�:"ᥑ�e������ /[|���dhdx��','�z4R�l�������e������/[|���dh�x��',' CdJ�H��OXN@�F��+)V�RNX���(����x*�NX���(����x*��NX��B#���0<a9�]���	�	��H�5OXN@�F���ax�r2D:�F���ax�r24R�l������ek�����/[����dh�x��',' C#���0<a9��G#ŚF�5�k"��F�5�k)�4R�i�X�H���b�(����x*4X'8a�,p�r<,�S��Oeq��	��T����,b',�SY�NX������Oe8a9��"p�r<�e{��Oey���Oey��	��T����,�]h�r<,��=8a�`�r< _�	��T�NX����@��,[�Є�x*�|',�SY��MX���|���Oe�/���x*�~ 4a9���
4a9�ʲ-MX����p�r<�E���� ���O /���x*�|',�SY�w�	��T�NX����@��,�/Є�x*��/Є�x*O��x�������w�w����	wy���]�a��]L���fw{��w�}���q |a3�Kù�}�\�d��͏9�^;����i����%��JvwP�״B4�pMKD�״A4mpMkDӺ�4�ߓ��<P��]��d#��T8��ҟ�Y�M_f��@�8$�(K$'��I(T���H�C`zs�8d��d�I��%h�5
f|	���C Uu|���p}W����яxr�O����R�dd��T[Hք!��&*��U�l������IU����F�ֺ'�K+[��z�V�������k)u�:R��u��yT�)u7�P����(����(�H]'Q3N u�Di��u)u8]'�R��u)u8]'�R��u)uU]w�n�J�Վ����2���^�4�w��d�^o�N�����l���Q�|��j�2���|�aV4!߁iYtC�L��P\��aZK@�ڟYȁRP�����т�<����.Pn0��-�P�x�c���<f�q�wH��V��k���LW`�U��պF]��@�Xt땓C����^�i�S����K,��E� M>���-ʚE�[��Tݤy}����.C�𼠶� [��Ā��h���/�h�F�h�F��h����H�c�o���瑭D�h����Ѷee�:�:Fա�+��CޑBnޠ��e�n������]~�����`N5]gu+�{u�7㘖+����2��>BҪ���?����54�_�i�S��J�LȞ�jp�͊Z����um�jә�i0XL��癹�0Xdm���E��8��݂���z5m�5p/�<�p
�y�*�����p�櫋��8܄�5��g�z��|�yt�����Ypvy�|}�>x�摽՛��Y��?*���4���\��/�kh��ɦ��"P��l� cw�����g`xm��(0M���(,�B�1���-��-�X�۳{���'PM���^y��o���v���J(թ�}>���aBU����_&��b��>S}��Ҩ��`��[��X�|k��g`��[��X�|3j�Ϡ��<�gP���j����owq��v�bM�n(�L���u�X��t�7�A5]9GF�A�֪X��<��k�=`��PM׶�`A�PMW�50:�����4C��4����*�-����ϗ��K�}��ޤ���n�����_�p"V����4����I���{��Ƭ3}�>_����=�e�뿿�K���M7���q�~�8m���q��� �� @o#@���F� �m�`�y �������H�{��<� s+<ߞ�#�� ���"�0��|DP��/���8�!>�!>���?���w=�!���M�g�.��@U-={��	/�q���"�2��ܲ�"��K�I��v����@�I�	�Xa�/�UFP����䯾LxY�u�2���껒AhL?f$��b��;kfRWo��=}Z�L��	@�C8��Gr& ��Aי >�3|�g�`� �1�� B?LQ|h<�@� ��	@��B��G�& ��A+� >d4|�h� ���.+{�Ćg	'M�˱��V�zԻr���| �Q �E$��GN���CW)
�^�N�������
��j8jWK��5���DE�@�k�����F01á���r�j�Ӏ�����DRM����z7=�nVnz�ݬ��@p�f�'��7+i@`0M5��CSq�vNg��M�A��l�A��� ��l�Cs� �l\�S�L`x�L93JL�A����G��ˊ�	ͦ1͇�O!�g*@+!#�ٌ�RI��?hyx�A"�h�x3�D0	r>�A�S?�s�P ���^xrP�	dR*N`r�J�%�f%w��@&��ssB�����҇Q��3Q�n��r��S���6���% O��+��6>�|�7��|�7��o �)�6�?���65��	�65��y�6�o���6�-�Y�6]Ġ��6]>�9�H@ SǑ`@f�#��M$G�O�6�����.G�	d��YF<G�9< dʹY ϒy� ��n3��Ѝ���n~���L4 �4X8y|���x �̀/}�+/��pf{N������yBE<$򼊯@N�^M!H���($�T���'[�`D��u�}�L�qa1b�s�ܬK�3����@�l&R��A����=���/��,��ϖ� >�)~�o��a`q 9��~
�:�\Y`�@! �
���/�Ѿֿ����!���f�Eګ���gI��y�&ϔJ�`��	 +o'����x�4˳�#�q}2)຿0:xA�Ї���/��5��� 2�F� f����b���>˓�H�ԐS	��9��������'P�K	2��ˊ�b��gȪN ���gY�9�� ���\��3�� ��7=���� �i�g<G6�Y ϒ�}Ʋ�Q@<��˖ݳd�'@�LO� �+� 2e<d�x<ly�<����	 �� @&��#�是����P�4�6��,���y?��#r�>ڒ�Ea	 ���$aWj�1���KBp~rz`z�� ��`	 ����e������ ����w����݇�x�_|����a8P����>^w��}�J 8��g;\�4���M"��C�@��qY�(�$�+��.�ɟjj (�eJP�ЄbO	ʖ�P�Ğ"�+A!�Y:<(_�B���xP��
�!������P��ā$�(`qT�9q ��%KX��,�@K��Pqkā$V��9R��.J�ΑzThwQ�w�\sĜ~��Mf�	�ļ���:fo5���"T�O����-�� z��)�����(�$���DA0��*��BX��[�* (4	>kFQ�I�y�	��(T-��EӘ���q��o�
���|���[
w�0�?�� йx����1�Ą�D�ќ"�}�H���4x���� �Œ@�i�|��A��%�����s8	<m+	�-�ϯb�8��$жx<?��@��9`/�>�������1?�wLI/_YE���1��.�O�� Ɨ�1�$1�h�	b||������G�O��;M�?M�?Z|��b�b����������� ��w������1>���������'���] �_ �->A�/�S��1BA�0�P��!wC��A�jO���FX>b�$�ѧa)�wB�0Q�%��B�PP#�'ϨixH�#,_�3�"9@�j����F���yH�#���(5��b��a>٥�!�C�PP#̧�����^1BA�0��S�ڋ!F(��� �<$?O!?P��b$����v[�
j��5��b��a�AB�Cj����F�o�P��O!F(��;�<��S�
j���5��b��a���i���8N��� ��R"q ��s��Jr�D1)~���<��LT�����T�� 1��'^/b�N�0W�/_�sLꉷۨ��� �;�|o�����fT'^$#_�dXK�����@q[y-���	��'J��E���+���U������B]��_K�x���@q�-�������j����Z�E���0VVV�V�VՌ$�╕K��/��g%9Lp����b��B��?����_�x��܄�W1lA�ʕ�f���ͨP��֫Y�0A���B�WJ~͇�ћ�M03�	g��:��� /
5����B�B#��i�����(/Q� ��,g�ƨ~Y� �	.K�1�q��. a��9+w� ���r���H�\
���ތ�
[�gLN�	-��q5����q�܂у;�0zX�W3����Y�A�]�&�:&	���Ò)"�O��L�&;*31�?����k��!�f�TfS TF�A�g�3L����9�F��j��'��0�13hn��/� ��Vj'k�Q
s[�Ь��ʃ�a�z�t��J�,���uF+�������J�,�����b�x�V�(K +��q-K(�V�ՄjFV�ր���a�&�Ɗ�ƚ+�z�x+�zB�Vv�`��r��r��r��rj�ݷj*-��A�*�F$��,
+Y�r�izф�;@�DnB�Wl*��}����Ml�TfX�yԪ��t�c�r˚&4�u�q��2��9����J�@�&6m*�I��rI�L�������]tA;��v@�g$shz�51�v�S}޶��bϤO�������A�g�Wf�aH�/;;�eεщ!�^7s��ϴ�]0Ѷs1�N!Y�c�+�/%7v�}P���u��1M0���]R-���w�wv�&vs��ϴ{���w�;n���_���u�x�w��T���L��u*UPi��L��fMp��VNh=��\���3�M���}RV&���R�oM�۹��A��kB�X�|���A��e��24�K�w!�g�o��<Ϛ��9#�J�cI�ž�C�:߫��A����i���DH�Xw�a1*΄�֨ԵN��?P�����Cb]��b�G24�e�7ڦ�l��s����?H���2��� �HϿH_Inf�&���d�`V��f'E7�,Pr(PR�	�bs�ԓ��a0e=(���dU`.sRts&0,=:N�&D:6t��ձS,���}R�|����j�!�&�U��!7w�R�Y8CZ�J䒮k�*�Đ,D�~����r�Yrs�>�~����������R�B/� szC�� tC�� �CyL�
�08�z0�7�r0;1\�@Iz�r 71g1�&�l0�4�w�$�Pށ�M�b��M�./8�w���Pށ�M�YL��	��l�6Jn[���h�2!&��tFr�9�Tn�HH�4\3�V<�O�^0&��݅d*�fv�R����������w:��OC�(\|��E�<.��y=ʋH֭Y!fi�"�e~ez�pQp�n!n�l�m������O�w��7,����=�����4vF�?<�;�S��?��`�����������ri�ٺ$?�k�K�د�.���{u�W�I�|�q,*��w3��5�a?����ނٯ���x���:H�&�0"�(��CdRǼ�ܤE���q�q��Ϲ���$�쐬OǓN������<�C�dt5>�"�XÓ��G��n�gM&zх�PR7}#�h�1�l��c�f��Pɦ�&��nh��d�>�.	��{7�m�p(�k�4�,��N�,�܌���8�Vd�@3�3���;i"1@ǌS'��v�dp^��J�����4�ÐIL3gh� R}l�C뽑� Uˌ�y�V�Dݲ&M)c�6t�9��TN�Z�$���]��%k��Ut�S}�J���`�s� �4Q��%�wm�ݡ�t��:���۴vvir{�%k�'��=�ދ�'w5iK���*1]�!)g�{�c{(	9k*'Q�9��g]np���Zf#�t��8�������d���dK��d��d���d��`[��d�t�[����&���2��+��Ɋ���Ɋ�m�Ɋ�z�"ġ����MMV���!v��8,�S�0Q�THf�ǃuz��g�twP�|�'W�:J�=o�\=/��u�	0saVM�Q0ս���9AsV���Kث��b`ď�7�� T|��������\#z3����-&����v�X5��L�v��3fB����e4.VY�����x�j.0�Y����M8&8؄�#�3���[*�X`eo�'�
�D����4�w��(fS��������̈́�&B��^�F�֕hd�c�G��0*���ތ��/�x��� �×�Ts&��V����'-���K�s	�2�l	��R��`<�	_@j�N/ҝѝ)	3(D�hJ5U�>Tj1����T�?p �Մ��U�
�h�u�����s]�@�j�#��9�q��T�xI�D����M&�]�J���{N���oB_2c�C�hj�xs�sOe�@bn���o�c��c�f`�Q`.�cn�c���l�q�E���R�j�4x#�2g����@C?bhj6 4p$�f�F�17Q'x�Qg��w��˘%ԡb��8�.g�u�X����_��Y$��{�%�� ����x_��������{�%��.������zGliV<��q�3��������H�H q@��~�a���'�h������Ŧ�o��џ��.~���,���x�$�O��,?��O��d>��~���O��-?��O���>��Sx��O��Q�C|bG�q�("�%Gıۢ�8rK��G���)��=Q�O�''�wd�(�)��%;�/���$'%_�/��<�E�|�G�Ȓ/��Y�E�'���c��D����%?Ց���:�E�|QG���/��wU�]}�\%�ԑ/��:�E�|QG���/��U�E��J��#_t�}�.���|�%_������>J��#_t�}�.���|�%_��/�I��w�vOvT�o��ݻ��y���]Z#�ld��FǢv�uC��;˽�wV���w��J]=m*�x�_�ݻ~�Ϙz��䳳FF�V�V�f���� �1]N�.w���>��������}�:N}R�YnvV?�9֊��fǄ�W��w �DۧE�NZ�u�YlO?� [-���؈E����|c�2*����>y����>����W_�ݾ�����@+	�����׷7��
��[�}�t鬺�����$��b�M���لh-��/ �����]���w!�'��͇�x�ꀞ�]^��]'���bϖ���}�?t�k�ݕy:&��	����i�������y,t��D!����Q2O(�%����Q�O(�
%�)=�{��	�c��/:�+�Tf����H~uJ��-O}�Ş�`?}�/ǡ�l��{Y�S����9��,����߻
���}�����������;Q�(��~Z����W�������>f��W<->�����7���R��w�7yS�&~��_//��}�?}���L(�w���:iǋ��������/�φ�����\�n���~w�����w}R�I�%%�}��8����]7�i�G,_��w����7PN&s!�(_)��:ѕ2���<y�z`IK:�5�aN��UC��*t%���XWv�?ܔ��Y9��2�;��Ӈ �?x^��e����Q�
�ULLc�.V �,V�.V�f�Xѷil�_�����������$��t�LA��r�� b�.�(� �P)�)�M���r��b�.�)���(L���t�LA1L���Y��F�T-WқD>Ao�\Io����˕�&Gw��t��ޤ�MЛ.Wқ�������dI�R��7�%&�M�+�M�	z��JzS�t�\Q�,�(�ߧex�,9�x�H~��?�#��s<7~B�ӯ>�}���=㬉s��������/����ퟮ���S��J?fO���?��~��~q�����f\汳�2���w����c{��F��>5�g���:�ǯOPL�y�����W���OR���Q12W�Rz����w����?��٪��+��
^Yg���>�+e��
i�S��n�&����,�X'�t��b�Q�d��al��"b,���6����o��٧a0&X�yp��K��U�=a��»��n�M�_��Y�6�1BY���\�˴^	k��>�*�;A��^�,���$|���;	�&�u֥?�u鵽
V�|s�z.Г%�M����,|��/�^zů�2�S�Ҥ_�$ |E���o��m>�R�7i�s�-�g�J��z�m�5v��{��Y��7��m>�,�W^븳Byk/�z%t�ӄ�B[�������h~�6�f�ˮ���y{�O)x�2h�E�~ES�o���|Y�P��W"�ʚ�Bò����I���9�6�}�UZp���1WFɐ� �;Ai^���m���g7ECv�?4j�*��z��PAJ���((C�+��_�{��o�𙧡�rF��H�'�0\:���)�V)�W�@�^�4����6ߦ�3[���ZdpN(�����f�'�P�����h�y���/������L�_�~���u�0s�����Mw���}yM g4�"�!WA;���KĕO�>��:�h���mB��t�5�K*��u����X @��pw�����2�5f��U�N|�J=y�*�t93zI)+��0jF���5�A����p���x�<Q���;z�Q)��X QK
*&a����Q�S���Y%��d�e��.��&R�doQlz��b�C_���؃ �&�,69-�b���(6=e�b�
�,��Z�D��J�I�T�Tue�I�Y��g�}Ϊ~��	q%MZx�ݷ��I��մs��'kX���"3�b�絒5\;&���h>»�J�9^����.aR�L���Ĥ�7?bՓor$���73
"a	����+���y���Ɇ;y��S��A=0̓�O�M�㝲������ҡb�q/�e21��i~�q���[��͍�����}ɲ]�
,���nc��CoE:-�\o�&9�R�+�M�%�Jx2��Du"v��+T����{ѵV�N@H&\H���X\��n��S��,�OgI����OF������i��z')�8������࢏]�T���C��s���e�ޜH:�h��c9��o��wc<	�C��D���͜}���a�}3i��+~%���[��~���C-n7$d���}�p~�����M�a߸�#J}R_�A�?�e����<-nJ��u��-��T��ɾ��I��ɉ}�b\��M�Ak��	Ǳ(�r4�DY�5���{;���bϤ�~���Y�{�\ٝ��d�p��}㓽�X=��q�I��IjX���Zz��z�q1��e�kB6z1��*)I��T�OJ&EI�	R�u+�s^+�&`�!(��yʐ�ӕ�(;���Ϧ�����0�d�F�� oO�� e�0�՘�^�LDi��A��R���]�U<}Ǹ���Q�W#�f]rmH�����'�1Cܣ���<���ϓ����������dH%�� ]��WɜϿ3"Y`\���ֻ(&��H�f�>��Cr��i������i���4ӾkX�{�z{g��m"���'�)�s>��qx�g����-������/���_�������_�e�ۣ2��*)�dR�$-y:��U�(�Z�eZ|���C�#����}�ҽ��SI��dEE�d$jք4��a��b�\ � ����G5�"b�y������Q<�ͭd0��c�d���G'����i��1GL�Б�Υ	��V���mB4����d�A�D%{�T6jrN�r��(�6�A>�l���RV
�m���S[U8�[X��;�o�D�!���U-S����^�X�"�漥_�J�~�ӛ,��dY_ii�N��������R`���J�	��2'9Q��!?Ƌ}+��u�����:�*���d�yퟒh[ND;	D&���;��;7�d�A�6&Q�m��:�|řP��Tx'Wl����v���&���-�KnxH��n.N���C29z���thb�Ti��}#��q�<O���<�vf �5^֗�c>շ��C����˼�	g������J+�龠?�N+qӵ�d���5]ױ|M���ڌ��E�lArς�D��}�KqH2���e7F�F*�ܵ�C�Y��_�uޤ�D�T��O�L���T5RYax��Xg�6Ҽ󬕍d�D�Rʖ3+��,9i#�Q�)��,7���ǵ*١;��F�,8A�M"I$R�S�'�<�{Q���г�X͆��I�X��Ɖh��u�	�}�H�kzo�˴jQ(���z����W~����$h''g�p<9 ��m�Y�P�Z�ɋ�dN'}W䠁�%�-�2���q��'���.��)uX�˓�oBD��Cu� Di|�$��?���7�G�DAﷶ&�а �N*�R��$5B��cCǓ�;ŢiҢ�'O�Ҵv�I�m�p����\�������Uб��_�����?~�\��~k8�?��^Ã�_���٧�{6.�����~��?�4��<��U��TJ�$f�Ι~hB(Nj��
�D*������:�!�H�C\p���L�?��=����>���ᛝ�h�+n.fޅW Y?��p����g���>�:��������b�}0,�\lQ�!'K�5]�b��UH�p�ްt���A�'?����a{x���R!rv퟈X�g�O-Wy�W����Qvg��I�XcYk�cB��z�8k
��H�mJ)9�V��!3��f�|��e���u�A����D	�E�r��T�l��ɨn�a���4��|%o���G����0�5iy{P4�
:�9�E�A�3(�$s�����O?�ߌ?~�^*�k���S*�n)�F)��6�~p�5>�%�I�L��j�¸���lT]c����&)�l�^%S���%?l�X~H�� �?�������n=�h�I�)���f�9-�L~�-g���H���m��Z$�DE��2,x۳!���^�i�Z%��Q4>��O�>�Ƴ�'Zk��Z+�W�^��&��q�Sa�ɦ�:�c�D�8��;��y'?�F��;�]���&�W$/['�)ٱ��67��\D��83΄��A2\N~��'��1��_ބ�RH���D<��vVV���iR�T$����}Ƥ���`����5ڬ+��a��s������1y�ڷ�o�������������˜v�&��_�p���{��seR��8����@�o����P��E忍�H�oc�]�}~�Ǯ��wݗw��������Oi�����&��ۻo.>���_� ����&�N������7������G���͕$��N��7�,)H���ؓ��?|E	-��7:t�o�o���i���o��xw���������t���������܏��N��E�%.��)����b���.��i��'�N�
M���o.~L�w*C��]G*C�N�$�R��ɐr��%�;tQ��شx4]���E'�X<�x��ă��cTL)Ш�i���a�)�C�	�r��!I���Z�p�FŪJA/���s�fǽ�d���|�UgE���E7t�t���ƺ4Yv�����?�c>6,��Q���Yr`OG�W�`T,T����ƀ�;�T_l�b�O�z�pa��	�&��Ę3�Jf���V9��IzbS���k���,�A�5*d�ة\�Jy^Qj���R�B��H�"�P�fC�2��ʐ(+7�]N�@��dJpc �7.w�ӊb�O�`jb��B��N;��봊d	�q�������e�r�6��B��c7M��,���(��)xʹҧK%����X]�^���4���G��H�UE��H���Y��`�� ��\��e�piq� !S�X���m0Vi�bZ�d
X��5y�\�TʍUZQ���HM�MŏV�y�V�+e@�7*���*KU�u�񶡖�}Ͱ��HbeH�Ue���B"�Xͨ��tX�V�ʑ�*��>�)�-����+�b�UE�LJGŜ����*JՖ6�5�ZZ�%��#:��bm%�;����Y�� ��v�©i+fa�e��'~ ��֪ VV�m���UE��;���Nkm�V�i�KY���<��-��qBŷ�>�V|�mT�_���t�
Z�b��nC�Y�Ҋb�O�@�d�e�+��Vݱ�H�� �+w�&�4��W���T����bU%I��\q��A9wF���O���g�����B�W'|�ٿ��c VT$g�5����b�N��e�����xBE��N��VT�픎Umo3��@Ây3�Z�V��h��-��V�h�R�-@�2.Vq��B��2�@m1;:բ6����Qw����)f+�ƪ�(���v�����o!�8X59P��6�Xż������!v��ƥ�����K~�<+w�\j����1v����B��h�nx�K}���ޱj�H� ��q(�I�i�������:.CG,w��Ն3�Etu��<VS5�ٜS�4�y]M�^����MŅ��q�*rpj�B���E���*�*^u��z	��r��+�����^��A-�5L��� �m�д�TZh5�c�����J$��C.X��2s��r����F�A�*�F�Y�yˢ���-罐�O�#<4+^���F���u�%OO�R��iNGX���R}أ3�z�v�KBb�T�,ld�~�AB1�~r�}N1�s1��C�X�u�y��|��c�r˚&4�u�q��2�~�t�,h�Q_�9�r�f��g��핡���Nv��e_-���Q��YFB1��7��i�h1�s�x�A�Vf�ؼ����cw��]��C�&}tL�B�h��.� ���ى�����������M�g��[���Ŝ>m��'�����b�C��_�����ֲ�������!7����N�:�#�:���B��'!P��`��s\0N�O���Y=�? z�*%j�ީ")�ն0�]0 ��9 ��u�Y'����N[F�Rٛ���ڕ��� ��8����d�������BaR�ʙ��NE�U�������cq�}�F���A�.Bq9��&�����h,.�M#f�Y�D��u$0���fn�\��f5Zڠ�H�y�ۧYhv����=.W�Om���Z��ƪ>�������jd�NrQVJ�o�S�(p9���B����V�u�րE�K�4ӭ/$+O^���ˇ�yʽ	;Ҁ$�%�-�G+�a7�*��4m0�ԣ���a���ڝC�c*H
p�q:�+�a��vX:��D����0CB�6��zƕ�i!�c!M2&�Ԡz��@?�>�`x�q�X�#� V>߇���!��v���~��	2V�Î{�Y��\,�b�q=�4��^�d��O|��V�~za��}W�v!��p�����t�a� ���_����_9�8d�^_�P~�i&����B�y��+�Y�ܵ�qH~�D���278�F��JR+_Q�Y�6����b8A���^1�+���p��AX�y2NF��s�ثu���U�D4��{�pt�G}���6�ŊQ
ǒ�\Im\�	��^y#mV�iSp׊�h��!Ј1�d��K��btk��y�b%��B�B��C���>��J=�H ��Η��^V0F;���.�S���^R0r��e��.���s9@{�+�o�4���.�.Ӛ!��*E,`~��*��F�H�<��4L���B���R�/�q�ӚUc����%��1��iՐKȂ3]�T0V��D0Vh�u�F"gj��aZ3�"@��R˂a��Q���0�5�iZ��iEZ�e���ǔ���+�Ю�F����/��B����q:�<� �8v%w	3�ū�ga#��.&����E�JX���C��rp>��6������#cZ���IG*-�&�T'�_L u6��?/��x.��|�'}-<�P'�.W�2%����܇+��R������(���j��4**yt�:y�.W��8%��<@f�����n[�ւ�b����lȻ��W�tÚ�5� ���ZQ�T��P���rB؊$��!�����,e[9`v�4Z+�5ب��<�'�2���ںu�ZNT"�j\*s��MO�Vo�*��Fk���B;t��ע0Y���Y6��_|q��΢��Ʋ	Β��g%s	� �b�Z��l��[�Fϸ��=x��HP���lRb�gQ�i�$�����7�;Ig��͓����͓q<^�1�c�y�K�R�N����3~������A۱�S�Q9[y�;�R;;f�J��U��f��F����2
8�O�����h��bZGa�n���x�@�ڝ�0�n\��R���x)yt/& +�=���J�aǻЂP����
�];V�{��#Tl���C�M�8�z)���:d<R���Q9]ٯ���>�r�,wB׀Bw��S0�X���.�
�v6���,Za�x\���j������Uە��ݳ�{�!�_:��.'d%���_��/&s+����\�Py�.�ئZ)q �祴��j� `[�E��D&" ?��Dd�g�P� 9
,V�����~���w񾿻��>\|�%��������ś���������C�ַ?^���PK   ��KU_�6�3� �� /   images/062f1f9c-d785-4821-8269-cd0e0f0d9a41.pngYw4�W3��(�/�w�X�{����%%F�]�"��b�jj����Z5*�v����QJ������;�w����{Ͻ�q^���;� ��9NCCDCs�@����A\���`�LC����}�������G���1���ҹ��*Hw�ռ��EmU���A��8��n�[gfQ�%�?�`�ҁSP�c1ʻ56�K1,���3B<#	|��h���"���H�w�vYv$���O�����ݧ��f�����ȝv�)�M[2��jS� �1T��#��2�AUXYպ����M�`X]����ƺ��z{����c=b)b?5�����u��d5V��n�J��E��B�"΍ p_� Q�`��8sD�v��#1B�"�<ӮÐ�>U  :�>s������(�;�]SM�R������QSQQᶀ��a!�M��sQ|QQ�e�`NB�AoU���&�Ų�b���\#���
,���2Db!i�8<��A��|S�%jsR<�]�ˊ��7w{{{y`�R\��	D���c"|���H{>4�8 ��*_jf�����aD֡=W���'��Rq2�+�	��X�rV��Iy�lJ$L`�r�*'R���˘1n��-���Hz{X6��f�a��ʩ�`w�#��A�������E�θ�q��`:b0��k{t���!���)'G\?��/��&E$����)
C`���ސO�_�>w��^��`A��$���	P�G�M��|01����7��)��EJ�<HdZn[��ú���+�J��E�7~�ȕ�v����w�C�3{���H���AӇ	�վy#C��TH�ɼ��u@�I<��8�@i,S�FIl���eaEfb�e�"x��h�t�9������:Jʪܪ��Yp9�9��+Ep���p��6��@	��|(N;%j�F1�G!ip�2uA��ʘ��\Wo�$�m2-���X**�(H��������8���𢃄��ٴb���Uᇬ��g.��s��`G�蒢blb"���!Q'3.K��[�ď'`᯷1b`�� -�j<(K&�ѫd��r%���ꉀ[��ߟ[[���G�~K.T�:E^`$�:�20�5 �;5�y�Hy��Ov�Â1GM��D��J!��h�6�&Ĵ��UE��@�a�ś`q�˄�h ���ϴ !(�^���&���SS���5�����g3Ep�5�qk�|b�ƪ	5�	�i%)��F���sF�]��ø0�i�Ts��ߝ�@	� ��-e�9d�no��͛�T�B�Z�	#v����2�tO3߀Y� ����eεV��D}�ʎ@b���K��xڀ��N8���3G��s�"`E�V��^Z�[s}�ǥ$�' �D#b���Y )1��K�RR�)`X���"�;��'IK�ڲ�ЇU�O;c�ꪐ�Q����e��K���Z.�I�ǙKԴ���4�Z�%�խ���I�0.	����
T57���X��p��Rn`}*$-��#5�5SM���hVpk�h�4����?������@+`A����Ҡ0�NC�E
�̚@x�Q�I�j�N~��(824d��K_Ֆa�.&���L츒K�ɵ y�!�Bw��~���э�3��D�k��+�6__��Ԍ�dP��)��z��LE��� ��c/\F��L<m����$�D�j��\eojyO�+�q9t�F��)G�}@&���`�Bw�˸!ʈ���<�$�ֱq4�/�]���qri]���&)C�>#�v����̼l鐗#X��Ch��Y̈́''DiO3fGʢX;�!�e㊺�LL*��m,*������+*���C���
�ۿ"D'Hσ�����t��ղ�w�$h���&Խ�j�ǄR"�M��Z}�֢ҫjZ�QY8o5��4P�$@�b(��r��O�11[�s�}��Md��X�K�P��|BC�h�`�c�K���;�y�.	�
O��l6��V��湙�&�Ʃ��Rmo.��^���!k�h���X��r�k���#��:�ܿQ%�n^iXA�����q2��RO��#��|���O�H�xKq��L�A}I~�0�u6@U%:Οz�&�����	�۩�:��p���ƴ�;��>�t�����Q7�뻳h�@�U���c0\�>���X��x������HҠ��V�vf����ˍwb*�*�)࡛=dg@k�@�J8�'�� ������r�jX�lIL�/Xxq<���&�t�zV㜖06����V]j��BB2��%����Ph��sȻ�1Aq���Z$Uph�>}�Ԕ,]t$��`�Cc�t�P_�a�2�m{*�[[�������Z�]��԰fq�U�T���B��>�C�����ҷ�]�U�q�[̅9�����F��!"�'�택{2����XL��,�g����ԭ��}4����-��X%q��zj�&��"}"���s� KT�>�cS�*�:�4M��.UR4qm�a�m퍡g5^xz�x�j����T�K��˥G��lkvq�7^��צ��X������?3�Ly�}E�#D�	�	�-(؂H�@ӌ�ѩX�N���	�bdeSj+�Ew��թۚX�#B�������Ş���Ԍhu���f��j���N���ɸ��ʈ"���"N%�`K��"��&�i�0�
,���o�M��������'`;Z1�+۟qχ�h�"��+*���h�i%�� �E^i�K�L^P�}��S�A	��=�֨��=�n��$��_G�I�ӯY��EC����@U��{0E�������T��p_	�+p��n��� l�槥q� G������R�oQ�Xݫ�4_�h����wG�ۯ�B��N��C��(@���a�6�(�M����J�m��YZh���$^���M��޵���n�dK�(;:B�A�]��d�l#ǋ��n9�nO��>�;��W�e��=~��;�@b�p:����:�D�4�@��%e[�,&郥SF��i����M���/!<q	� q'0��f��K��Ai�"���<]�؃���%�����Gk�`N|���?��LS�v^��)���~�0�k���!fv�p�5̉G�C�=�T�k�\s/N��dѬ��C�k7���|)�^g��ZR%8"��[���q���]?ϣ_Lj@����ZX��d���ѓ}0�6��#�������N^�+�5�N��zD��|�h��ZV27w8-lBDt�)P�;*X�=@}ȳ<�i������ǽ�������6�A��A%��
z��vd������`Y_};��Xmu���ʋR/Wy��|"��-xuyy(�����ܶU^��4|q�������j_����,�t�>򏹧�TZ�*��dG(e�&#�.�0<b��[R|��p���h�-$3��
/�1'�f�Ԗ Z�`B*DZ��IUE�W��Qx�%�m a5O�(��+3�k��Bh>X78��d=c9M|��~x\T�A̦����1J�����"�������9,�|���Kw�of���;fw���qo�M��4h�fZ�pI&��4L�Fd�^�wf�"���PC�:��ƙY%��i���׭0��6l *���OJ�f�!�#�����t��J	Yz��F:���Z^��M�g���0t3��j��W��<-�.��Z��Xrs�_?��֖�i�l��5�`p[Zu�<�.n�ۋ�S�U-7i~�S�HN@{om0������t�Gd�<	cA�efXet��`|���\���.!9���Rǰ�\����a�Vg�Ry��շ��q�����s&�rí�ȑm��P��y�z��� �P�����U�b�eɫf���8X1�	�ZwO(6\��w�����$Jb�{�|��:���w�M�c��j;n<�@27Bv�	�
J����~wH�a5����Ž<���0x�̈́�����f&
\���`��yz��꾠�����`�#ψD|���n���"��>�\,��o�q���Zl@�i��de��UL]�D���|ꟹ�8�zO1��~)�����)"�6���a���\�G{W��9��&amK�;;�҇DCa�q�"�
��� �0E�=��<���r�C���+��_��.WV�7{h��ץ�ĦE���&k����#�rY��.	ngP]���?38��ec_`�*I�q���(��^�g]�P�3{�� Ax�+��?'Ц2��&X���0��8�
w�&C�?p�?
�k�@�\�#�I4�*���K�w3i�1�򘎀m=�Y9�T��ђ�oM�q�����PCd�q�Y@ʧn�� 1>�`�*�R�6�P1�(2R�T0�����|�`MTH�����K��1țY�fV�5Ҟ�x��p��%"NH��eF��ڣ�V�T��ʟ�AydNu�Vrr��"� �鿄j')m���+�_�	\p,x�c�'ʽ6���.Sl#�b����{P~�Z���[ mK����1)�2�PR���wbgj^0� sC8�rt���2I�h.=V{s)���Z-\�2��>���t���-F��g�z�
���ʴ�7F8��R�r=����[�A�ģ�V���V"c�"��rؔ��y.[$�9DM
�Y	�	������DL��^&7�oe�A���L�Fh�qP��#����$�"�}w���p�)i��Ł�U[�]R�%�q?��ɓ#����Ū�ԛ�j�Ҩ�	$�N��^�!�����B#L�6γd��=�چz+�4�ma��հ?ʥWa�������-v�5��jOs���X�uUyA�����}����z����]�f�1\!�y����Q��%s/�o�R� >�/�t�~k@*��4��
����? �2�VڠfH�v�����S���|M����I<�r%�xف��������RM�JYC׃A9E�в������>M��FP����Jx���]p�I�F��L��-�K���K�S����k�^��������3��)�fv���	�h��Գg;w`����|q���	�{�����Y��@&�J�U'�'�F;�/��`Ě���Hf����p�O9�)��{����S��a.�;��ۘpm�!=��@y:NB���OqA�����Ե�k��ȑ�0SKS�2WX�����P&dK�N��aWظ<h�q���x���߭!��2Ç]L�H��Y�7�=;d�\���2vP8�l����"�� sh(�8T��:Y��/z>���@i�(���4*�{�K��bb4�	��l7�WIb��|���*������,[a�����Uq������&̛��堟�]ܾ=���Iq�j��0(�Օ�� �B�EL��!�T]��A���r$�짉,uIL�-6���ZS�@�T|^����k0=ϝ��fl*1`���0�/�hj����v��-*�����PT'��F8�M��/������y��sOvFl�~p1�d[�:Mڑb�U��'h�GDe��s�����TTW�����cR�D��\��i��yh��||�)�v������Vj��!��i�G�%�_D�JK��=��t�)p�?P��R5��r��*IN��3�[�h���K�����s��v�;%<ޮO^v����TJ�i����o Ȫ�ȝ�0fC*˒�(��qb������������h6K�!�.=�R
%U�ֺft��D�̼�zrY-�(|�JJ���4�8�̞<Q|�ell_�c����jSI=fZ��kAԲ${��Z�M����t�5�Q�438�䫩$��}���b��V&����TS�C�I�����8���2��'����V�M.M�I�j��N2�%��L���NU���#�g�_1"(�}mT�������Ɏ���ۍK~w�� �&kJ!�#J=�UH�ǃB�Pn�]���¢'F&<^x� f-�����h��fe�J����m2�)��0��W�ڴ����4ֲ�\#*��e(w8���a���oI��{��Y1�w�ұr��΋�x������X�jh#빢��	��E�$�`�Ю|>�o�@xǨ���òs��%����iA�"/�h�]L����8�V��_o^���	�d�٥�n&�_����i��ލ�nW�$2�#�iT��L@�z���Jq�.Bt��7�'�J*�����A�s�h�A+nP���,W`=}=S+�_Z`|���5&���W4�ʔ!�^�w�T*2QX%&zY
b�`Q2R>�z`l�j[�M�	d���X�\��O�j=��^�i���9�w�i�L��jS\�;�y����Ew�hM7�e��{x4&����ޔ����N�Ƒéc��-�*�����lSNi�g�����)������>��%�ej|����!y�<�*CH����-5dĒ�=�&'t�.rU�����ˑH�]�Қ���%�H��� ����V��^Eæ�t���G<(N}HV!ӈ���摪�w��%Q1����C�2U])�,o�Ɖ�p*n���>*n
9��_л ���F��{JV]�\�0��))5qH��M����r:���q�.�HX�(F���婦Fx�jm8mD�i��g�[D��jT)�B�������5D�ߕ����� 7�`d�po~������}C�]Dgm�ѿB$k�3��{�;GC
#�ks���b+R�X���O����u#�n�?kG>��$R� �s�UWV�C�0���w_����X�����ӟW<4e��6#� �W���oŅ�,YLZ�=��X#�}�4���e������m�X���I}?S����Q��JGYд����P��pו+�x��)�7�u*�W�ʲ$W�-|s��z��qg�w:ȹ ߪ�M�4�\��������sM���l����7�4�Em��͡���<����-n��QM�j'�5&P���w.`<�� �܇�}�����G	��oSjS�#����ւK�����]�p��^i��8��i��T��0��~��v���FE�o��SM�ޮ�X/�dv��U6ɣO�XZu�"��5V�=;�.x��v5����2`���TȮ�*���/�M�0K��%;F��f�� `����VIk9�������_w.lD�lS�;���׍�^'<1���$�m���s�˒�~�]��K�܌���۪M�/��I�	��.���?/�Rx�L�lݞ[�l9:���ԡ�H=w,�Mɍ�5Zo<��y��RQ�vR���iB�l�x|�gwo�����v�ǩ^�?4��06�M:,�Σ�z����s�ٱ�E���[���z-U(|M�-߅=�5������pٛ�?��q��~Y(
4 :�uk�r��#�u�u:�A��>·�IM�x�����C�5vi�-?�*��g�7+q��Gҵ�u� ���ڻ����m�r���<=��Z
\ҜCq ���j��@�LA�����
C	���P��+�vD��]�����]�A�z��O�l��_���.����Y��n׬�b�=UX��a�dD�@�a{8��ʖ�h����J��-j�9N�k�L�4N�$'gkjG�?nX8?���:�ǋV���]��YfsCGG�A$��kG�"��m���M�Y��w�U7}G��e�[WC�"��5M��lS�u�ﾪ2�i�{�x�T�<��d/fZ�R�pD�c%�kx��3Q�j�`��t�!���/wm��ך�E���w.�^�h1:���ve�}���c�������V1VC9ԧ�~�i�x�)8��y|��g�K�&�%<X�HRC��@X����ߋ�pKXo�����~*���Sݫ9��S�G��Jr���D7�]de�?6_�*�+E�E�	�{�n��Y�%}\���fٷ�č��:x���d':x�"�"�f��?X%����鷀��]��E2�&�~2~V 1���8Č�Ļz��^D��}	�4�Y���ߧ�1gjO��&T�,.p��d��7�ې�5�N?�[��~J6�ܨ�#FP�xX�w}�2�<�!l}�d�G{}���6f�&lA>���f��~X����:�Y6���uPr�|Q�V�*�Z;瑟��'0�'���翹��ww���[h�o%�}nGٗ��
�U�o1\yF����GR�񺰑��_$Gp�/+��<�]��M��p�uG����;�!�"�C���t���M�6#7?���_^�}$�ba�p07i���;���;}�S��=�"��`$��H����5n��g8��7�N��F���Vy$�c��'�"�I�ʛ�����!�S�j�D�m~�]X��7x�g�L9����=S�^>�b�����{cxi�G�\p�~����&�����'�L�q�m_��4��`��V�{�`�[Q+��T;��'��V�"�ma����ޘ�m��쏭FF���G���|B�ͽ,�`3�%H�[uI��E�d�P�J�A�0���kJ�b�]�~���߇v�3r{� '��TZ�\Dl�N�Mc��+L  K�ƣ�b"#��g��~�]ڦ��
��������*��`��9룿,Y+,����Ye�n׹�0�2?��X�/J�tK�,���ԋ��7N�s�e���8xܾr\������q�+k�Y�g�e�|�w���޸�X�Y,+��r��Mv�����>�.��ӏ��ݡ��U���;��q�2�m,�fk�#�J<9�άW��c�Mq\��9r�0'�#�`�[]��Iu`��/
�ŋ�����rn�B���|��)���j���]��k��{����\-�5�$��bܳ��{��?%Lۋ�3�e�u7�2���]�ak�xY�^x%�M�$�=l_� �����}�ë�90���<����0P88!av}jg��^�
�E��߂_�<-kU���E�-�Ųf>��'��,#�#�ڞ(� ��v�U��}y�{z^a��ʕ����}�J]
=��ͳc�{�϶�*N%Ɗ�y���2�˵O/���Q�hf�z� Z��2��,�~p^�?�h�%ѯ��,��WU�������a8V�s`�n�E���9�ߺ�_���k�G��u6h%�g����ئ�HR��q/ �����f��h{xZ�7�hh���^~��#£iô��_~s�G߄�|_�l����j�6sl��#
��BL�~l3����+�n���ڿ�������'��V�ܜ��K���y���n7��;v%9ow>i�tߏf��q0b-Q��Q��M,h�XPU�v���vg�׮칂��qɰ�{yG���B�`P�L�Kg�.��		xNzu�"���j���uN��������a������{�]�lR��G�\3�3|��s�����|�F�:/|���5����\ֲ�ѕ���E�S����ݪ1�{i�)˚���Z­�6;�o�-���gc�����p�n��Y|9����ԅ�X��<\�u��vKJ���p�#9qF��2}���-��>8�44�]$)ڼ-`�m������� ¾�$'�C�3R^�����g��P�]���Ɓ�������p�/��}h<��[��������ՖX������^���͚��M��TU���_7��qv�X�\YE���s?A��PE���j�yQ����F�����K����&ů�0�c:�g+b�S�o�y��@�=
����>y�X�(�h�P�]�U(��{�yi�7�=}˪���U�Wѣ�Q����1�/L%>Wļ�B9�$�a�CU�{�X ��l�l���HΚ�#����� ���p���+��}ۇD�N���'����P�6���PQ(z���Ӛ���^�s�҅8I<�JѿK/����_�d��Xi�%v4�7��7�	������2��fg���y�Z���6X������V�~�zI��E7|�"��0�]-V��Ծ�Lă���Fh��㦝��PWRl՗���֒R�����_k�2��yԦ?LH�l������!]�3*��y�1%�[u@ߝ$�$'�i
����Ub��g��(��--���v�գ�����0������Mj�]J�qx�E�/���3+�����H �-�>���E�曛7~�sr&'���+,n��e����k�}����{�Y5*Y`����pKftz���D�mB�|�He��k����RXZ�Փa��L2ժ"��cQ���Y;��;�y��O�SM��	z�N����[XQ"6q����җ2bᐒ1��a��ƻ�m{:;~�ѯ#���ƿ���:W����i��+�3�Hl�jk����SU�Yת�7���kͻ�w�Vz���_��{_,��Sm��C�`���j'韟]nF�K����� ����j�2)w�z�� ���:B���[^���S�=���΅i��>c����s��AŅ�M�k�o٥�Z��j����p�*�?��뮋߃��>붙���i߱M�V����W���K�T-bڛ�Bv6Kv#�y����.V�K�858<{�.��������s��0����y�ë/~~<H��]���mq
�Ҍ�):���A�h��w�{��%��ZjO>���R�6Q����vO����V5D+|�Ga���-��s���[�rJ��f�Ei0b�X�o2�ڋӋ��O���������$���g1E�&��ؤk&}OYo�W�Vm��Y`�L7ɞ��d0��lu��B�ֵ��a\\�w�n��w��i}�5ո��O'�����+M~ʮdY�g�`�U�A����	�m"������5PQ�"l�i'�G/N���݇<�`��=
8�'�-wZ6��i��q͍��;�����w��9���~o�ߑ�2��&�qw���)�<�%���,*_��ʕR�P㰃'Eq�����4�ub�'� ��x��i�����t�ĥ���בb��4�N鲰9 '��d1j��P�S|��x4?6|;�	��[���R���r�u_��u1���(�t���Ȓ#Y^W�A���)��"�1���p׽� �+C���_�S��˳>�X�x��m�G8|�=�3S�<��t��N�<��TH�K#,j_�|��a�^���{��$���)���}��-��ΡA����ب��D�Ѳ��c��d�,���!l�0�֥����ȋ����?;/w.b��.}���S�GT����ӻs�5wB�3w�i���~�Q���XV��#�ߋ�������S��t��	�;�U�h��uO���-d����-���/�ݟ!J�%��cb�yD���������Y��	��+�KF-kb����dq��(��T�ճ��杇�=`�B��(a6��oT1M���\"O2X�/I)@�m���VZ�&�8�6Y��ʖm/Q�0*R��ly���0K�|cY�����ܢfx��������f`�CsPմ\�nz@1.��Z3Ƨ�`�f��m���{n�H���枝cb+�$%3̘r�U|#��[��&�32ejw�	�ʙ�\$`�3LI�j�%\4�0����;{S����Q������W��C����ygP��6���veW��vq��$1��rk�]��O᫏��ϗ^�`}� .�@�;~[[�E�yUd(o����tZ����,��Z�pf��5~���)�4����k���4N�|ع�^���벃�b�����h,�v�^�K�˃�pYH_�b�ߝ�K+�P!�9u�M|�u�sоG�����mU�nq�r�����im�>63u��oP��#��ZA]��w������?�ٌJt��)�e�S�t�:���t}k����?�(��P�!�P­��󜝉���o�����ͽ����r�c�(���dI�(��@�A��+�*8�!�)V21��ð/�=�=^MQ /�����e(��N.��Fq��H����-��Пh��'��X��_\�� �pl�do�{\��y��_�+~�Ο��Y�6�p+�y�B��f�k��`���@9�1�#�,i2�u)w0s�|"��G��}s�2�~�R���{Ik��\��K�+�e��*|�naS�C�A�e����+���Bn�����=%�^#��)��qn��&�3���J&N�E�t{�	���9-�	|.f���������I����_m/���L*�6(/n#+���ʉ�F����8۹>�]pL/s�!��ר*�,���]���N��*.��M�(��z����ݹ��]�n�����͋#o�=.`9�vYl{ѣt���̈́-�?~�j���>x�wqJ�!��XT�sV�w��p��2&�R��H�_�E|�0�岫��1���#w�jؔl��١�����]�������io\���ؑ��Z��R_�w�A�?�9�������<�;����%R���oB��M|]��߾}S�}n9[I�
9N�ք޹w��ʼ����v���<;O̧�Z2ŗ�ٶ�e�t������p0�)wx�P�������p�^�Hq��k:iTY�ߴ���On�ڏy&7�FqJ�bt�3盛.z���}��v�f�\�����(�Q����]
O�?a���o�9�1�����g�m��Ir�j�́iH"3q�<�R+E�*솎�62��	��+��]�o���zv�H����*�p��3���=e���$�>������+b�vӱ��t�o��w��t�ѭ�ם�f<�ڭ|!C�'x����C	�2Iv��	}"��-V-\oq�10��ilƿ��C8XjsC�"o&����tL�o��V<�!yR1�2T����Ų6�s ��_[�X%�[�Uߜ��.���Tí�#�O��� ����f׻ċUR=ܢ�ߡ8٢`�����TAT����Q��w�d��Ʈ���H�o�!��Z��;_҅���}�pb�6������5����/�9H�\*Q�'	�~^��o��|�͏��ewct��Q:Oj�H'�]���Ņ��=J>g.�dI�|&~M_�������X��3�&4�z��=�Ɂ�2��v@ٚ�����~�U����&䁶m�-�:����%�9=��S�j?�y��m�
���BY/>���c�%J��C�n�t�A-J9JM�T�
Pu�)r��n#�{֦(9Uv��2��1��l�D5��F�)�+w��ۈg)j����h��0	��?�|���h<��;7%�}��a9M��f�tﯬD�'K��y��A"A��Pr��?��t�[xD�f������n��\�$h���J`}y��곻�=�O����,�<����ׂL*2���i��9�J�'Di�X;rpz�}�K�M�ܡm@K8�kjj� ��(ad�5Q����ȟ������͚�¥z��*'�t�"��������~�݇�>:�4`��x��:E��ۖ�'����C���{���T]�cn���䲱�">�O���TV�`�S5_�`��B�p����Q܏gC,K�95Gw���$VyFj�z���
'�n��w��s���̺�#����%
bP����7f�5�����c�K��md��WƜ��V*���}���)�~��pY�5�:8���������������Y0����e+�Z�4%B�1�	Ϲ72�b���
��_� ��J�CI�˟ �k�#��0��C�S�nQ�-�c��@�3�l�J8�l��|���Pu`Y����^L��]O��q%�7���6���~pX��W8�"�C$u���͵��%$�q�ւ��nm?I�x��D��Ii�xz�UHH�2G[����؄�&�W�(3�'�N�����M�&�/�>���UP\��-T�I33K��w)��Aw�<�wr9��p��\��=v����&�����Ɛ�,�fAN� ��RJ�V#8���h�@�&kiz*Υے��1Q_Ҧ$�R j�ߒ.���|t���E�eGDN�M��5�(y�8$J�F��|]�����;��}�΅��iY�%�ūҭ��آй�=&���K�LY�隹���(2��pR�ͧ_�6/?��	�z�����u�?�0�:.S��%�x���Ϟ���/��hR;r2�.�
{f�ǫ�[y�����7��}�E*"�I��N������7�Eu։{������ ��0�ք�X4(�b3ע�ҁ�}6�Ϥn�U�º�ϙ�~Yaz_my&Af���p�4��.���>e��~��C:̎��&�H{��Y^�A�ӂ-�%A˓�7��F�������E��"��J�Q�f��R۽J�$Fw����(�n�@�7��H�����c�z��PE�*�@Q�@�����dD6���M�Q�-1w���K �K��0�wݰ�����OW�$������Ô�HM5�j�ݿ����<��T�����(?t%R�-d����6y����wq=ڠ�x#��Rr�le�|��,�#0y���OjGےw��ot$,1yk�,��4��s�@ώ�UUЗw/
&��ު��Xs���Rʧo>|�Q�3ϋ�N�"�Ԯ6�U0XG��C�Z��ݭ���z��I����D�j�������r/.�ua��#F��Wn;v��e̩f����ߥ-�J?����X�r��ؙ��}%�`;"�!���ҝ^xi�dc�oa���e�Ť-�>��_t9%�X�qW�c��v�t>��-Bڲ�Z:�8��3`�O:zȪ,����[W�j"o�I��������[��S^�~�;p9z�~OI�_��Mٝ;�A���s���#g�ی��ۿ�u��^��{$~������˃��n�>i� =�=k7 ؤ�I,=a��?{��k\�{�ML�R�t8��c�W�O5��տ~�r1U��=����-����~��������ژBZ;2�?��kq�!%�T~Y��O�Q���Y"���?�:-�w�;3J���r��������8XNV�iK���D��Ȋ� ��~��+L7O�e���1X�j{tgx~[>VY��ڽ~�x�����l�Њ>!�s��k#��6�i�uׄ��y�e~��J;*7տ�����`������F X;ݕ�rm� �5�����@�*��<���G�c��tFkqK��jҏǍ��p�n^@DD�%���)��2��\\v��^�H�X�֛��oۧ��	-Ӝt���λ$�ο���X�վ��W�p��m-���̊��Q����� �W����w�R���$y�2�P��fX^��h9n!�3�y/{!��]�}�#J�)�W����鍏O�t\��]��Ol��,V��w[�$ߝ$h����	Ԇ����Q�/�{㈁��-:�N�0/��n�%�ڒ��h�]B����\TNgn��|�M]�}��m�X�ٔWl��:�}/g�� _'��P�.v�5����c�B��QO
��\�;]I�Bc��E�gd�
�Z����3e�ˡ}β��H:76��s���*r>����b��Gr����bM��3m�*�HP]�Eqx�v�(o��y��ؗxWq��~��m�}����C3��nBm�w+�u��UZ��i�oi��$��ı�ی3ϻ�2I��&��d��I��J�6@c�'vg��B��L�������g���ؑ�E>�j�x_�|�R�c=�ې,'��������]V���վ�4��A��"B2�<���/�V�%�M�?�~ӹb�������׋�����5Z�ܹ���`��f����UxK�?^)����~�9�ۓ��σ�����J�͝�@�^�|>����t�m,�{��U�c��~��y2�|� +�	��nSGڠ��K.�p1cqB��8���n\n�k+�<u�iغ��k۝�j9����
���l�mk_� ��A�V����ʋW�@	�S�"��Tt�~�u}�õ�P�9��IU�I�>[N��bۭ�d�4�����{��_��E�y������H*O�<:�
�������m��_>������|�'��-�+W���N�>�+$u>"C�e��V>�EG�'�ƍ��!K�z;Z��������,_�ٺ.�Ae���F���h3��O�"�=��U�_�8�N������}ҏ����3L���=3q���e�g�U��7��-��#���8��O�Jk�����Ux�G�$ކ����ht�d�h�#]���L��n�+�$��/�C����uBD��@~�W=�]<����^�|�����Q�t���x��8Ϻ���{���oH�l-��,�I�7,�*pz�L(҂�
�g��h'�R�ֈh!qsUB�Q�X�U$�t��kiE�o��Yj���]O�-E@Qϴd�C���YGE��A�K\��U�A:�;$AAj�N�QJ�Aji$��WXJ�R�%Db���Zj?~��qϹ��=s��}�sf��e6V]�!3O�������	����TT��71��v��(]U�g�1FLJ����֟����m�q ��U�1>[�l=<����6P�������L�cXk�\�5s�;픡��M}�A��������7��j��}�Ԭ ��,fÖ)�D��k�:9RLc��%�o�z��.EeTJ����ϒ��{|f��B��b��$�t���chO��oȷ&���Zf������wZ�.}Q��)���nb����'w�z�%�����[_VF�����	�W�D^J��	
��!v
K�i9]
��yܝ[���������ޒ����Rn��gj� 	��+�
�A��»:x16��~Sf�&�1�Ł�l�Ԇ5
^�=�	�vhA��i%�&J�%�Uxң��w��T_럇n&L��|+��T��³��&�E�<a��3k��ip��FMk�.wI3����0��K�Zgz�����sQ%�UNq�j��� j��2�\GD'b�����i�l�)��O��I���
|&�o��h�N��;8\_���=�,2x�����pl��dMG�d�����6�%x�91���A��vt�"��Ih�~������T�a4#��#6:�{�H�ָg��_��P�ňy���h�T�~ҵ�ziڕ����dP��g�����E
���\�?���!>�;4|u&�8���P�v0i|[M_R�yb��7�Ai���$���.�/��X}�d���Vpm�%p܉�������D\O},|/$���a�u k/G���e⫛�@S�<��j͊�ę�o9�Oٍ���-��0?k�̚����@x�$�]!�YQ��Mq}��˦�c&7ʇ���[{ge/;�%��Y�IF�����7&�1��l�"kR����t���[Au��팛'v�0� �1��v�Xu7�6��
Fq�ߚR� Y�wQ�_�kF��e�f�8d�z��\�[�X��^}ᵛ|] �f��m��z˫��������p�^�Bz\��F�I�0�o�%GlxIvv���q��\�۴w�g8%��xd�<YN[�-���p����B+@�h��F�&tf�����$�h���+Rc,2A~����[~2��g��E3��PU����X����v��H��h����,��6z9�8��J���߉0�Vn��*&s&�'=��FzVh� ;�R��C��r�f�J�?��H�T��p[YY�Ԛ��:�<�g�-g�I��=4S5���{����˗t E^��^sɰ��@_�R�y�I�E(E�������>%���͂zN����(��m)���K,��ￍ�Y��ή��j���E@�+�>n�gJ��.J����mq���بL�\���^8uL��}T�%��^:�Bٲ�F؋S�D������x*
1k�X�/�5�4ߌH����{|d;n�r�M�Z0G���6:���JNE�I�B�ge�d�%$'"D`?����7�<m4�%yB�%��������r @뉶�������+Uh��B�����U�;��z�y�BN%���5�Ls�Q�T�`s1�Jc�	s]��	�-*f�IJ=���]Ɲ��������X�=6��)r��El�>8�	�>?���mъ�����+�p�0Sɗ6V6��C�S��s=����G����W翛�Qm2`=�٘U���{r���Qc~Gq��>��03�Җ.Y�?�B���ӹ�m ǹ��!�t+��q������2���4ߓڧ�vOx4X-�F^�w�w����j�s�֍�n��d�������e�/���W�ns JD*shHs�NX۠+,���Z$Z�T�<Z�s)&��m./��W�mlF~�|m�����S�~�>��D�mR��bDi�D���w:���#AY�ɑ�ߙQWhT��x��� 򔟒rT�t[�4زuҜ�fV�Li�
�����x�k��/K���JK�����x83+�~���2{.vp�>�K�S��~p`3����n�������ٕ����"2�F�R��;��'�$9��C5˧=��j�*���z������2�V��]WE��ۢ�pK���Y�"?���"܂i�p�������$��Rx0��=���$�x�
&�Rs�O���	}���+]ʨ���i���Z�P��܆�)J6\"^P�u��E���Θs�8��F�HݥJR#�,�D4���۸a#j�/����,g�������Wqq����ri*�2q>9��7A�����0�$ 2ΚYejZ�)�x�'�m1"��t=�OƄ������*�{w�	��(�XCJ���F�����8������O�P*��:
��y��4ĩ:U�l�9;)���]�.��6S&*y���^dÒˣt��$y���רb������_�T��!������"�/��c�$vT���c[�h�K���O�Q�",���yF��1�o����{b�4��~�Q�ɩJ"��Z�WG+�������'{�A0}d���������a��hs�f�=٘���z���;��=�+��BUM܂L�{��7�����-�	��}��;��������ҙh�0���s��h��>�v��T��^ى��_au�|�<V|e���x�c𞭱�<h���[K�(�=E�5�<�v��Fp����U�6���(z*��׽Q�gS���
M~=���pV������/��i�ۜz��(կ�7 �}��X�%;���'_%�ќ��LS�~�u霈��-����\N�b�$�ߤ���0���m~����t�ټ<ۇ�Ը�QIDl] ^s��U@{����/\�f���7��fz����ki�y�Zp5eu���`�Y(����6�qA��0`�����T���њ�CS��+�ۀ�݊�\0��WE�	��z-�>���ڨk�P.� �h �E�;_��9�����8)�%��\X#�/�`)R�|�`bY;Yا�$R"�F@�)��;0��>����l���t������v�]��^,���8� �
sI���0���n�>[���2ѫ�ܲ��ҙ� U}-Rp���̑��9Mu���p�`cJ/d>M�e;��%=�����X�Y�T�b����ٶ��3�|z�n�P+�Ar�~��uLs�=ÆL�DU}�`%�-g�f�����ވT�ՐFy�[�f蓜�a-,�p��vY��˘��M��Nܪ?ٽJ4��r�r�' ���I�`�y��eN�%z�8s����x�Y��Ϟ�ŀ�/��J�TT_�%�+$��[�1�*�.W*c���o��ß	\S�"PYXM2nA���N�Zp�]RFZ�=�O��6S��>��X��wUs[��M;B��{�2�so��+�:��t�m��I�w�4�l�h��}��Zh:,�%���_{V���R�Eյ}���3�D�8!+ �7C�J��c(����(4d���1 9�/���Q�|���b��k���o#P�m0.�,��N��o��t�t�����4����?�Ӗ�S�w<�Wm��96�NJ�_]ZR��X�샞�Gy9��b��9�,�x�*�W���p�W�8C�r'��7U�����D{��=z�6�f������2�9�8ễEo�iP��;�$�����-�o����H�"46++ڝ�_ϳ?鹞<E�싷#9M�|�':}[��\:jm�ߏ��"3 �侕�{W�7SE����5D�3���@G�G�X穰��Z�X��< �!�h���xw��g���F�T>�miЩ!IU�*����#�����I[Mu|=}Ϫ
o���O�%�H�=��N�������&�tO��v��ަ��lܷ`u�~�*�\5U��k@�*��gV�V�8tI�u\5pc�h'#�����K~{�Q���-��f� �k'���'��@+KJ����L�n��1�~R]��S?)!�I����i�n�!x������+�M����\�+}�pu�2q��?����Z]��o��\M�n��2��$oOl�DS\�#���yMR(Մ3��K��Z]��Ηo���;)N�zqpܡ"����TH��W���$���`���]].�(&�_TK^�6��b؋�'���T����L�+n�ڐ[Y���/�f��ZN{����K�Z��r�;���q��ʊIR驮�|r@�pc�l��P���`�vf�ܯ��g}&�7ҁ��w�gIa2ԋ?�����ߍ��� H�*����{a�տ�'���kٰ�a�$�x�iX�X}�G�(h����s��T�����l{N`e.�\��	���;�w���셎ͮ��i"r�[��3��#��$�o�Lz��6�E�7���w\~�!�|c詘I���u,z��l(�����Ut���O-v���\��/�ڳ	�G�{;l�?y(�Żd��_��95��*v�ї�a��Q���{�ηV���O)"S���K�V���Ф4�Hp`��6��̷�����2p���=�~WV.�vP�E%!������i��VC�Y�rU4�fs���뻹��à�lr��IBr:��S;�uIR
��ivr�2��T���E�>����ڦ2W�T�Yb���9�执Վ��Ai�׸;sl�tؖ�\�<���Wo�S~1�yX��lڻsǯ�PD?�ؼ�Ț���y���\F1�&�$z�"��;���p3_�@����z�A��T��6�9�Ks@r���jB2T��b�`�铀֥�h4�l�9c|�'󞣚�R3�YC]M�n���v�죭P�b�t��Qz�������J�~>�I��C�f����W�;V��i��V;'� ��l���G�(�1DIi�4唯�q��߼f��V^�;xuS!m�<L�t����P���X�������7Q� �w./:\�R5Oև!�ۢ�����|�_����f�5��M�@�2K9ʋ�D��Ź�J}j-,D_�殞� #��pd��u��u65���bγY$?:Lŧ�ȝf�&��e�`���֕�L��#�a%���ہŚF꽹O��ߘE��:��S����D ��>�~sM����C��g��e���㕏U�"ꐇ�����X�����y���~�zR�D7�F�2�J�L�͕ċ�V��Nw��L��L�Y(�����_���:�w�%�

���״��4��Y�� ��t���i���2fE�����3�kD��z�Y�n�q�|����g��j����q�J���8/ CH�����c�Ӑ��+���\'�Z��Q���Q�]֎�hX��X��b���=��ȳ�H%�����]ny�|u0xѸ
챧��&P����Л@�M ��Dy�D�⽾��R'O)���xx%a#���j�Uv7�#���{�n�NO{%����?�1�iL��U\�6�$�΍埿�wf�c[��lm̚q''�A�����1P�c\]Z�SI��}	�( P2�8��0��n+Z��>E�֭u7p#1Nue&�/5˿�3��ARO�u�O�P��6��o[�xj�Yd�y#��O"��애����V��>���ڿ˂״�^]2�0�����鬕7k�����?t��/}=��*Df��Ӹ���E6�u:���TX O{�M	�!�H��L�
��/]�M�S�HE%�5=��5�v´:S���-(�n�%hLn%�\G���b�M2��qEY�N.��Y�"�&���2=�}4�3{Y�y�)�N�	���#��Y��ן���0D�<껴Q�{�4���\� ��Hs=k��	�0E�{
l/�:�E���	�O'�|:Y���[�&�;�>�Jkp���w -��&NLB�k�8������;-�^�T�e���>z�G7��]��z�0��S��[y��E�?ᱩ���7�ǚ-���lv��-=�ޡCFIoK���M�9�Wߡ1$��(г��~�FA-ocgŻ���T}I�
�ll�P���iN���MQ2�`�L�0�5'�}�i9���*ahRakٌ\׆�n�p������Bk�:�b�HC5�d��y��Q��(�uCP�U��&vͲ��D����p�hüW�����n��3B3��ݠ6M]]�q�7󰛛��KXW`�' E���O��ƕ~	��n����h��Q*����Q���U�-�[��~���7�Ն��)En�����
�*h�&
��-���e�W(A��1+��,~�����/�L�XBoR�~�����[�=L�R=p���FY����aA����>���S��+���ge6(���g%nÖb�r["�ŧY�/����������S��@�v��TǓ��ܙ��X����h�N�L�����@"_�U�7h��86L�G����^y��#��́���ߤ�)n-��t�f� /O�˨��IG�*&`��kݰ�&�g��>�g};��o]�TǼ��yu���-�z�#cnҌ�"��������/�Ȁx�����im��i;�I��B�)��.?�����B=�%�Et%�7����#�Tqwa�z�W�.X)��݉������R�+�<��_�����	�C�bΒi[S}VOHd����#���.��R��Y3�*;-�7�d4;�����d}���Oz��B�Z���g���eW��UB��GH""�l��mZÅ?���HG����ݭ{/��'n�!���<�99Y�M�'���ޟ?�V����\�,�f0_�zo#<�6�bA	l��U�qi7|��m��.ߴ�f�>Y��0������wX��
k��@[�P���0V�7S61�����1�eN��3��@Y�;=�	�ga��m���!{�aPq�q�Jc��tꞦ���@U�ݼ�gk��2R�䌔�3@~)�����+���{7S��6v����1���,]3�����1�d��I�����՚���A[�+��_틋��;Y��'�H:�t\�c�����`���P)ЗSz����WS����誺Ow��r�ܤ Q���al���q�e�R)�ٷT����Mد:^����n���.��E�}�n�!)v1=5���̞���{Z7}��d�R�A���v�^�b����?@�YM�}�F��ث��)�m2�2w�;3��Y�B�Yh)rJՏT�S�D#���{Ot��c�]`3D�P�`Z_c��BxY�=�丣�4�_��ElCv����١lgH]�䅚�,�Xn?0@��͠�Zck)�v�>W�BD�1��_>ǔ��Z���e�e�G������e�J;V7�Z��9t��uR��Oޚ�jTi~����#�!@1�ʟ�5�(��;;��Z	�D��17�3
{0�?��2��0YMO�nL��Ia�/-�t����W}!흤�2��C� �7hY<��u�h��,��,7�W��x�P��M7��k�MƊ6u�4%��P3�� o�B�GY��j�.��X6v����s ��{�1�8�8��'�[T��=����$��z����O�c��[5q91B�ޞ\E'L�Ny�FtB��`�;`6e��q}�`S�|�	�8	���`/���-�J�)�6-��d���S��B܀#d3��ų�=�ldE"??;����>1�)��v.z�g@'7�[��N-L"��b��r�ƪD곆ef�b������3�ԣ���A£��������ܟ�RHn����H��G�UB����}_�l��ew\����O�^l����������JM=�L����g;]�#�^���}�GTX����ً��uk�����[��Z4Ҵf�՝F�_�vg��'�ե04��(ߨ	����U��B�og2aד�j�{/;���dE����+�%��k���5G	=������{��MԷߢ�.D`	t�AM�Ŷ�����������=/���=��-�Ȁ.���``!�E׫��� � �/��kx��x��`Ԍ~�_.t��aESxXJk��tT�jVc�(��U���h9��`��$�[����b�]�q��v}\�!BU���h�ǍHf��ܳ_qW#����l(�b"�`��'72����x$[Y�����9*CZJ;ɳ���w�Ml"[�U���RP���0\7>���)��Z-C�o�j��C�t�y%�/�G;>���zR�Z��9��rN������w\�8*'V�� ��a���y�\�d��0F���Ij��FO@q�*��֠Wq�9�6d�+3��k\m��E>d*���3�-)�3�@eYG7�]F�c��w��_�~G�$7����.�\�~�#r�
�R=�/Ew;`nCs"z������i�?�6bO=�[􇤖�'V�d��A^�S%�᪩'S���!�m.55fdd��ɷ꿕��pU��/�M��u\���5}D�e^���>��P�)x�4��`=w�����S�F�h���|�xssz9��9�XA�G_m�f��X�_�Y]�,^��o��/���(���|7;���1<a1�3�Z��%%v`�GT��޾v�Ư�йRO^~q��$�@�J3Ú=H�_�-�ﲄ��u��2�h�K,�����_���k�N���+"�?��[�)��q�:�]��\��x�w�S*�^�R:��E���q���&�+�7�[�:uj�xJ�P����N眢��%�����{v�AZ����;]��������ԮG��/��X7�m��C�yG�_�wH��p8/�^����0c)��{�:S��h�E%?�7�Y��^R
��i�U��r}�xm�5Q�?��y����LJ(�!T��%9��h
m��;�[�ǘ!O;;@�5���� *�"���矸���Z�7|J)B���F'�O�έ�`����Ua�����h���bA���nװas���Q!f~�=�&�B*���z��Σ�JJ��ǆ�JM�r�F��1m5�����x+<�şkiK����o��w}�_��8�=v3�Z��w���,��@ �1�C�6�%~k��ަ��ʋ��xr�jB���u
��ӄ�\�fPf1�"�Q ������}�����<�O vj����©�A�Ͱ��[:iF��fN���z����6�
.��e����v�)���[�W�X�FХnKGf�崆������w�^	�,�=�@A�M�+qm�+��EX�5[�g�#�l�_�on��3��M�@�U�
�����3�d���s?�9��և۱����DsF# `V1S�տ�J�"{O@C�X�熥�8����I|J3�����ޖw66�l�|r�w�Ӓ$Ϲ>RsgX~�jvA��Gڌ�=rj�B����F[��ysj�<2���O�FmX���"|�I�dbq��Q�X,��r�k	Id���gJp>��dF$%WR(.�~d "%��sⶣ��Sp?&�E=�]y佥������6Fr&3d��	2�66��.8����錷3d��X�(��E��� j)�	S�y����D"�!�e[����Mgv}:GPa��e%�`�b"�.�����6�W����'�h���o�~)�iiYf��+M�Ow�`�o#y�o(�̽�*��h��x�v&�T�[��`��zǪ��<�����$Z�ͯi�l��̫�H�nJ�/���n�y��k�uipA�.�;�xYB���',�m��KROS�tn��20�h�op�M8�i�rt2��dK��1)�iG`�����{�Q�/�Z�{;�w&�P�)�%� 73��� z������W�?N�|���a��8+�~�����n��g����e�s8^,��r9 �)�����K��&U��R�>|/Ȗ�V�!!x0��8�<=�_��DPA.�w�Ś����	z��p
833oq��
���NG�"cL6��I�mV���O6��ϸ��@���{s����)+���8D[��)=�4 !	L�����FI�D��iJ�c��y�^�Ub^���꽎9i��v@�د��ޖ�RZ��Y�0�M!*��-XDҢ]��R��������a\��ǞJ;���4٩�@�:�60o"�3��_�������ZS�h�^��<�<�J<�[Ԫ�dd��͈��߱S5����kK<�g�8�w�`�Ƥ�yq��8v^(��E����nfm �p�z�6���O��JR��n.0�W���SI��K�	
cd��7?�GM�C�����`�=ۿ�p���u�0�����t	���W�<	t�>�*�qĘ?��c��A֬w�~�Ɓ���1��E6ɮZU[�b5~�l�z�%��|����7`���������#
�`�L(�lȫ#a��z_��߁����k��֩m	F2�=o��}�_ܹ�*Uފ�����)g�&���W|����\j��<+�:}e\����J;����f*�d�Ό��Ɏ蔾Wk�x�
}-�7$��^�c�bs�_���K���xr�X��L�|*t�ίz�`�k\؆�cۧp��Ww;b
9�_NO���V��ȿ�F_�a{x�:mVh�'�,��D����Թ�[`�
��D���R�A��kp�7%����[��8�S���{���`��g���b[-���X���M��s���ٶ����G�4=XN�N�kd^T�+��&ݞ��r��=�����@U`ԗ�b�)f���!�j�7J/�z�̵/~^*���4��ɥ";l�ن�-���Y]9�e��ɂ��q8�g�H����'����?ʖ/��kP_�^�/��7;���	�ރ�ؔ�z�KD�R۰5��V9�+�F�I�xڝ�6�@������\��\��/��U���k�G��"N�`��~��*}�֪�5qp��u�(�ɘZD���(}��4����k1ƨk���=�����VPc2��A��H����K.��sV�!�[��A=�ʖ��=���,~�q�
�,�d���{K��X��D0�H�K+=ܱ5+��J����?Q���#�ǫ�}�[d�xa����+3�GgGWǂ�\���)F5b�i��ڱx�_9}m�ln��w��d��݃��{�1��!�&��ĩ<{��4U�ܫ���41�����1�VmǵfM�ZIR�;�,u��`n������\ox���7�6aO�3��=ZA2AW�	���]�j�y�p���/�������'�}��&��j���eV�v�g ��#���e2�����^����h\�#������t�U�}�Cߪ˷�eRj�b�L�M��v%��^M!��:<�_���B�J�S!���
�Ś�W#��{��M��oe2_R�u��'����թަ�{{̎h���*�f���lҒ��e�3(���l���H`��{�~rBGr�*���zlK�y�C�����i�#ʄXUu3'a��+!�u韆\Z�R|H�&��|1�_	[_E�R�\A��������#���F��M��5��x�|�^>W�͊L�����%O~x`������f(��J���LwH:���{�t[m��S��SQ�r~ꄺ���ixi�R�.�cv��F�����q�O-������nBe6r�����la���ZLC������Q����ش��7!��2
y�����h���~�D;;cx��}��d���n��r��v1=c�քn���N;L�dOKwX���:}4|�C�	iE�[�T;ˎ�=_�������t�㝟a�	ʣ�8<�zӡ�◇ffw�zQb�$��=C��&0��ۖ	s�ڝJ�����VM��"��Gf0�c���y��7�y�������3e���*.�uS����pn3;�(��Qޭ�u��V8�V�9��)��	OHH�����+�7���f���G�% �qA�!�������IK�NU�M�|��H˙� ��`1
s�/�*��g���7�y�`<�]�`T�ꊟ8�&¦΃j�b��ji�$p��|/���z�C��r��vBy�,
���x9��P�?�[;�sC�/��n��W�P�
��T�T�ԹF����D;#���]�gR�[�[t�
2,�#�5+�i5}�
��"��J�M��=�i?IKW̛�j���\�z﬊����u/}�Xt�ժ�̑[�y;�>i�$+�B�i'�����d@��]��# �o9���������u�^*WF��!���8?��rsu�E��!�e��?������}�x���=�=����)��ַȦ�sg��.ب�|�V�p���l�j~��>Z���+Ԫ��eX?��&�B���4�r-�� �?��5MG튎5�܈��Ӹ������z��"���I�}����!�����U@��#����C�Ft�Bę�>*��(�6�,\UzM�,lf�������[Dp��ed�;�RP�1��&t�}Z�6�n7
�@|� �Z�G��t����c�M�m|r�4���V�2�7Z��-gN�$�����mI>�P����uw�w�����卿�]�6�mmt�ܐ�T�'�n)�΄nk��X2���a}u6-�O5��u_���q�sQ���J5ż�?�C{�K�z���u&��'�_)�c�3|c�I�L)%�����d���^�܌R�`F���_?]�- �d��nT�|��7k݉���LJ��?�*.#�߹7@;Y�^g���Xްf�oES �9/A�z>gB�ݧx�^��~�����5���>�  '2
�!��V���ִ�LԮ��F�"6i���cR�j��p�d�j��{'�+�g˧���`�T���H�Q��re�9��A<�ay�����z(T>�\����S[�纻�~4�7|>B�d��4�lh$6w������f$H�̠N����!�h�[.E�+�,���g�[ٙt�|�����T!���A^�C�P��\3��z�1����O=��JiF#;G��m�p]���^mxI��VB����W07�C�=��]��b���E�^Q�1Fu;ųV�t.5{7��d��1)�M?�k�Vdh��?A�m����岳�.p�H�m#>��a{�kF��Y����3���ޑ`���G�d�6BPNi����p:^,�(h{�R��se�O@Nt���CO
d�/���4%i��lsʟh�5k&1��A�,�М�p��nF<�?H�F �C�V�s�;5���^؜�e�%[�1٫��C��x�h4B<N�w�F��o9Q�Zs��du�Z���?�9}��(u�@�Y����x���L�cޛ+�X�Rݣ��B��_?�f)9<,{S�XP�ې����:HIո[�U=B��@��Hw��D��~���q�	�q<y��nh��j|QT_�P����2��i��i��?#4GDH+ʵ*
���?��0z�֧(���/^pG�Q�*-)ѯ�������d��������.P���#а�I����Wm�F~9"�ZV�,Mթ<�?&i�˨��\`��3a���k]6&�%j�a멨޼��f�H��J͋�K�%{�)ڐ�ncO-�(|px�{��,���\��D��Aiٴ����rAw�F����	W�0�,y��peS�3J�HT�h�0�A��Zً#�\C]�ȂBF| f9����K��0~�EE�z���7VSk���@6pg ׽$��K�2�z#@pg�泤K���:՗�Ƨ$�E��bkʬ�2p��0[S��"
nzzJ�ї���8�B�h?BHf[��z�X��Lz�/I���P��U�J��fg�5�+�"{�����V��K��
gG��w��!��N	Y�����#�{��<�>og�ԒV,q0�W�B'���W�+�^~#�
�3��0�^q۬ 8�}=��8�xﱜ�L~���������"1'O_�?%��)�J�a��j��j�;H�98��Tଖ�s��V%i�*�ս�NC.���̣�Z�1�i�5	��a~`g-��Ƌ� _E�DO���F�Qql��������-�ϗЏp�(�3���z�|�`����5Cfkj� G9F��X�Ȃ�k�K������;ڹ1�s��g�D�ӈ�Z?��j"��h]����J��`~ÉR>L|lf�@VZV�`��z�x��,T���Z܍�{��m�Y�~�~�����1a
 ��'���#���k�aM�Iw����q�sf�*�V��L��=��3����ѥND�1����s�f�V�vg8gUM!OI�	O��`zB�A����\��	�����6!,�W0L]3��!�*y��Q*���s+���K�+�x� �����Vk,�,c1��_�.����/!WN�k=8~�ξ� �����-m����9�$�Q����aj�f����5��@�w;��ܚ$�7#2�2��5�8\6hW��Y�YB/�O|��
�G�F���c��4�M�U�s?���������PL��ڟ{B�g1�N�ږ9��~q}dMzr�z�s[���}⤐��-�O�ԟ�$r��')zL�ixʹ�h��F�2���P_���vn�4ƕ��1�˝��k�"c9�`9�O�pc��^���L�����G�V��,���^����	7|�e��LӪ6^�$�˂wy�c*�����k�F,g�[���xkB�j�2ʴ�����m�\�:{�|/��n�.*���Zͦ��w�A�#+�0ٜ��f�.z�d2|}�pM�H�C��9������K�Z�DΫ/���^w�I�i^�AY'_{c���>謿��rN�}�X�hk�%V�{േ���t���;XA ����C���I�ԃ>�ͻ���wy����jñ�ܱ(o����������=�����$y %�O�8�^"�,k?�3�]��X���3��)>�S��n�k<s������ �4��Э��� 0�I*�ؙ�����:�O���;T�Y�U��h�E�&��`��m'�"@�CRc��C_�ǶWWt��}O��r �)�Yz�n?�N��
xuf�0�tiMje#ӫ�6|�L]�)d�n��,������	��<8�~VE��|8�AF*<��I�O����o����N�1��[�D�P˺D���C��g?g՟\�Ӵ~fr-U���ľ��Ƃ�13����Ҧ�����a��-�x�L)����=���x�ޫ�}�y{�	��[/
���:�)%�h{:��6�����8�p�J��� ���,�!�����X�on�B�\�;a%��؀�O-�lb�e>m|-���֡1`w������O�\�=�i��%c|���&�];�4�|4��~k�q�>���d�"�gK^�	��%n�C���1��8�DN�^��;:!_<�N��� ��ܕƍ�=X*�é�f�m����X�j$Э���1�[WG�ƽH��p
�O0E0|�SPV7�m}�Κ�a��k�u�-�lHx��hӠ"�z#�֨�0���b_e(r�Ɨ�A �/��$�O����=q�}�P��TUP)����-���XK�����y��V�zZ�_h.`,�fnΒd�F�5�>�0�\J��Raa�
=�;g���^�ܕ����82�4C�<@ И��T�*O�<� ���t��;?5V+>�=�w��<͊�����Y��Rz�o5O�����6�<�|?���CϠ��Ϫ�'77[�"4EW�*x�_��1�_�qo�����K��t��ZSb�m}��!\��Þ����m��}�d��IK y���I�.g� %v��D�����㫋��v��d�����=���=a�8�����\_�kj�;v�Q^�8����g�+��R��������=d�E�I �ш\�Z�%_�m紙���a� �ɦ�"D_=�=e��%�7������.��wM$s�p��~�~:�B�=-!�|?S������,����EoX���fK��4���"x���j�Ꮾ�?�f���&��Z�N+���O󑕟@�����m�ٔ�ss�'��O!|�o�R�w�M^�+��as�P�պk�z��*�������K+s��y�3T[._�v"��  jo�x��O7C�I:��BBh��h�Ԩ�9����kdU�`��5����质C{�U4?R�,�� f�;V�h�f�1�҈Z$�����"��幄�/�cs=�O�S�*��1H�:.+�"��ig�1����㙜�*7��f�z�U0v�n���|ߤ��3<�����/ϛ�b�=�_�({����<��ȷvv�dp�R~hN����C�y!5�5,���L�*�����
D�̼���k�)CD�Ԕ�x��L �]"�����l�y����EQ����z����P;}����c��r
c3�qV�jax���fj���⬵]�&!�M�-���K�Q��0'p�5B�h�3��Yȭ�4�̔|�Xٯ'��Ȧ3p�"]�W"ІLX�h��	y���mJ��|�����p0�@�6���@5�k���:�=�}ܗ���BMS���5�t:�>~�p8�Q���xQ�EWN��#l57��7�<��)�dFh9RS�MSJ�Á�D�X�	�/��!��un��Tm�фF=:wRN�j¹�:H*49�~���~��v�MU7��l�l�����<M��r~8��=N�T�h�s��X��kc��0�o۲,�o��?~��������'}�v""�)#FҼ[)����4�D䵮���tDGrc��m������?�я����ٟ���O���0�$���z�I9��ٲ�9�|mtLIY��\�T[k��ə�sd7�CJ��5��F��)�q��u���[0�߽{/yZ���VuK�㯞���?�߿�����~���ǿ[���?�ß���}x�2���������?�/�����������g���I��Ĕ�Hj��nW���A	�8��s��=�����r�V�v�k���α����N�h�L/���r����__�o�ջ.#ڷ�c���a�kڵ0C ^��v��_[4ܛx��ķ����1~�q�qr݉R����󋙶��Pʄ�h*�L��Z]�j�I�]d`L��<M��pp���v�^�����z��#�Yۊx/�o$:	�y���� }��c�ҕ^�q�4w�t�1s�T�_$~l��mp�@.��,����|�]�iz||<�N�4����mi��e�-���~��u�,Sak��u=��h�Fc&u���F6i|ASW)
���]n|#�';�=�n$B��!�(��C��˺.�����AՏ��Sv8u"Ҁ�E����/�)u�bFDe.�����/�/�۪U��P��Ur.e���8w(���ű�#�����4�T���F���u=�'�`��sJ�X�Η�__��̉~�㻿�ջ�����:�k"�x���P�^�����/��ۗץ�)e��u��(�������0���G���iuӺ��b|Ş&��^^_���4M�<=>>j�1s���C�!�����CP��Xb
+ȸH1؉�o��v���z�]q="2OszƷ@e�i_!�䤿>[���/̖��m��Z�:M�t]n�ff�+,!h�p�֥	o7]�������>~��烶�\7�v;e���<�9S�,Dj�t� ���$��0DĂ����t8�R��TaP��Q���tտ髛@�a��X�*"�:d�d�)�ݜػ���v[��|�,�������w ��V�i��X��twoښ*�'Jc/������z]��Z�IJӔ��)�R�z���G7 3H����cXmb#t�9A)�J����C���k!O%k���m]kk� �a[���L�յ.���\O������� "M���i"�D�Y)��o��%�����?�o�b	�8<��u���HA�ޑ'0;�_���v=Y�	s���WO�_|���Χ��޻I��.�4Ω�v�Fs~8ez���.��o_V�Ô$q�N@�fM��)��,|0z�D2�sJP��l�{�������Oحe����,χ�}����������]�������w��ǿ���s=��<?�r�<���������w�g�Ӭ�l �j�\.O��E�M�"R�N]�~gz�&�F��� �,a(_E\���(�h�F<�d���ܖ�����[��С&��џ(�%"��Lі�m�=�9��C42�������a�2'&�^��X>P
"�S�st*���HR���">fwg�����P�e�-�u���R&�2��\z�˲.�c`���,��%��+��{Q�G��"�Y@��81H�L-"�sP�}��ǊmL�m mrH����!��T
���sj������g��{�����r�^.����I�y}4A�6Bu��������3�p�8@�(oa:�& 	�x��OV>/v���O�,�M��n�Pڑ,<ur�	fb(�=??�����O���p��ّ��Vk1��Zy|oO ��
�)Af��V��z����e]܈Y$I������{*v'��x�����������V
"�D��,e��a�9���|�>��w�?�x�����~����w�N3���^��jJ����ۿ�����o~��'���_]�F�Y�m'W3g����kl�Hi0*=E�(�u�b�R�9�����mѵ�˺���L󄩆�T ���� ]>f%�b�֋-�qƉMm����c��hܑ$@�RJc���7��s�������@�=���䩔y6�Z����ea��5}��!Tu3��l�뺮��)g�.�e��k�F���n�:��ڴO�,�4�3����u=�ψ)����C���|��f$�x1Bg�D���i��M��8o3�$�y� A]U�t�����@����md*��.�ryyy~����O��SB"��01doDb��tզ��"��O3�u5���j�����TRI������2�^�
r/pܻc���8�#��1���{�ɑc�S�v< �'�U���z�����1{/���R՜Qo��e]���������w���t<�S�ޮS)�����_?=?1����_��|���}E;%���w�k�+�mݷ��j]U[�ə�)���E����⧏�g��wN�����^_��F�<MIh��}���������������|zD��8�y����z�]IhLj3#o�K���-���͔%� wN�8�Z�۲�S�#�)�~p:��������[�����/���\���>�˧���7�|�����������W^�|xP�����
��L)�;�Bf󭘥�^�o�8�4�_�΂t�ȟ�N�$�ɖ��/������s�EP¤������y�(��T@J�x!�"����t��ܭ���YO�ŉ���GD��+�Cȸu��]��R��['"�l�h,M�n�j�7�uYS�c��<ϒR)��U��dN1�RJI�u}}=???��r��'���x%B�~@�%�"�,㯐s�����,=���-L�t����m"�DRD��0.[SfI)qw�tzyy����w��}�]�$:8�&�K��j˲<?=��_�]��p��:�l��`�H�ذ��D�@�^{N�̅�0��Ɵ�H��"g&��a�DC3sa��jMh�8��>�N_}������x$�Z��k����&������z��������n7Sm!��9��g(����'K(�A������Z I�<5wwZ�u�����J[>̷z�����^-�|8�ß��d��_}�r]��o��������?8�4��;������MhfGCit}�������	�W'��q4���f��~z�^[�M���QX�C�ٖ�v�]��i~8�O�4OeJ"N�H�0*ay�=Usw�Wrbaq�.����z�^�`�)�̆U$��SL���x@���'���x�̿~��!PLw,�ù��9�ᄪ����w�������Z{}}=̇�������xD^���n��ڀ=|�TK�)�i�
F/�.��KgT甧S�R�͒3'bauo���3ӗ���u�X�A�?8���A@*����X�4oa�v쪭���ry�����;�4�Ge�L�����ܵ��H��\J1���|���H�1s���\RNFlNL^[��u�q6��):r��e�0��:J��� ��O��ԇ�HĜ(Q&ml
�K�$��e]�������w�Sl�19�55������?~b�֪����:�P`��Z��_3��*�� ��@�������9Ȼ����a(�o����������w�W���>��o��L/�}W�K-%?�����O�������Ng:}PΙB�҅o���;�/f���S�(��� �f����"��Zm/�/��q�f��s>=�u}�Տn�ÿ��?��?��O~��w����J������Ͽ���s��МZme:�Y�,�����rE@�Z#fqg�3����?��G���Yix�^F%�Q�p�R����������w��eh�T�cRSbw�_L�Rf��r�Ze�$�����}�G䴍�13�$��pkfJD �����s��Q�D�[��UU�$�9y�Z_J	�Gf_j{9�^�r�%�<͇9�t��@7r�,�O3��_[��/�OOOO�?9y�j����T�%��!LB �z2�)�!������]��?��a�;GD����q(�H�M��f�'߽ *H�Y����������Ox�r��Z�:l��G��˺>??=?=�k�� '�$NNF \r�����1�i_����}/QO���������ٗ}X�d���$oX��b�IF�O*�u�m]�[[�c90����eYT�iø���,�$|ں���mYnU��v���l�s�R�$(ѠMgH�Ƿ��w�ڰ�G,"���Z�eY�C��ND����կ.O����k��|}�����?���A�ry?M�)������M�����:��a"&5G5���s�x����ƛ��Y�	��E%�t<��v�]�����pg�z��˫^o��a>N�y��������H��wN�U�ն�����f���2� 'HD��RJ��$a��DϞ�y��!`�i���۷˲mz&"�_��wTk%aI%����n�\�y$L��� �_�%��ח�?�{��x8�i&w�F� '�R�Bz�	�������|>�~��t�\SJ�C��S��α�T�aDF�����F{y{)�������3�T �B
Dy����K&V�Z����|�<����y�y�u"�?��r����zA_��MSɥ$�\&3'�p/�Ol��}�񘚇�
�3�1r�t#Mr�����b�.�|��F6��l\J�������Zk� *�sY�!vא�"Ԃ�Z|��)%3�\.�>c���޷ڦy�ʔK��^�F+񦴁����j��vt �#�O�;9�28Oڼf��E�������g��?������ok��Zk���e�������ש<|b��\�X �C�^.��4�h9ϩ0�63sf��ĭ�V[.YM�Z��������i�s����)g#?���ֵ�?�����;�Z��9��.Fb�Rr2������|��{E[ ����vOk�jK9���c������2���Pp��13`��PJ��#%���E��SJQ�NBN9�<��Da6�QL������}�V��R�EP��>M���ej�o�%C�7��TLМ�2]��0f��N��q��ג��k]������GS�$yU"�5�9إ�D,��R:'r��nݩ���< 	���Y�u:,�UN�D�!�ߙ�"i��	��"�N�Fe���͗uM)���~���~{8O���x�%1��w�弞�/�Ϸe�z �m�YG� PG����O��{�A�g0)c�PE]��fG �9��v�0�$�s)`��Z��R�䥨jk�������x:�{��t<ƴ�3>�,j�[����uYnF�ԅz�!,ipLK/y#���o�,�݌E㎶|��
���Ԕ�̗eQm8��fI�x�n�^��w�����wx����ӧ#qaV�oտ�n���������qK�(��0mM�C*;���%���>/
��ou7��;Û2���@�^P}tJ)�d]���v9_rz>����)F�K*��!�'��VD벞/g7/S9>�#œ�h�0M�jޔ��]Q{�(K)l�n��J�wc���_|���DP�Y����|���T&3[ʴ�˺,�5�>`[l���h�k}���������������áL9�6]ֵ����r9L3��n������z~}��һ���4C�2��S��S���	<4��1�&�4�7�pǞ�����z�h��y*E�RJ�a63�co��6m�<�
��QO��\�u�]������+&qL��J�I9�B�v�uY*�t�=O)Oe*���U��%1�d�ts&G�MLq��2�	��1|¬�<�T��"��2F�����������i�~	�8�г,�JD-j��&��o'b�眒 �`���v<DҲܘ1p���4M����XJ�����yg�g���g��`�u{L�f�,���z8��4[�d<yN߿��G�'�z��O���p��<�R�O���/�����ky�<���
Q'R�o���r���2U�);�,Q=��y�_�p��e�D�~���9�w��Oy"t���;�C�#���UkdJ���qr���)IN9R�L�����?�}�&)�a>OpW%�Bau��0p��;Q�\ɍ(�\JΥ0&q·9ϥ�df˺��)0���(뀗\�-8�'bk�!#������9��sLW��.�K��?���8�=��7f����z"�PK��u�`8�����^����|9ߖ��̳iUL�D���.�Kk�����;7O9�Ff���-����4���'�_?G��dNwAN�#��l�Fac����r&w#�+�ĝ8�D
vBO�'�������eY�e1m��KMRe�-6k�A7�����	�v�~��!���+�G�仛����\�9��׿zF'��m�'�vHtCaY\�ڵAP˜\+������^.��m9��>}:9��X_�����H���,�ܬ��0�\R)�ʑ�t2�]�8���ls"�QP����~ �J��\k���,�Ռɦ���Ǘ������k����w}8̇�������ϗ��֫ύg�obO��i�8-n��t��}��1�/HV4\�?��=r��:�s&"�sRJ�c`�L����N�j�p ��W���ݻw��)�"53��6m�5�":d���0��4OPu��	����1���_�$��n��S���T㹻�$!7R��J�S�,�K�����a���a�'�wG�~>�������w�ߕRN��Z�ڂ�xQm�>??�����<OXB<"2��VIb�n��<֐b�Y�B9���<���o t�>@�v�e͙�܈��12���1I�y4���ʔRY�u��#$ �������v)�f˲ 1ᇔ'!�`���Z�ۺֵA�ODR��@�\�ND.�nZ-$���{5S�䛛a&5NrJ������"it"hp�P�-%�%s�R�������� c`A[k����>,�C<.g&n�ik9�s)圳��$�N)�D_��^�UR�t-q4l��w�H4 ~�Sy���n�`���^����X��t8pb&������O^/�����sJ)����L�wǏ�Xy��$�T�d�t]�������bFnL.9O9e�6���쮭��Rb"����l�K'���o����?|��s&�I�9Jٝ\�4��K&��XDH$S�,iIy�懇�֚��eܔS��û�w��#����׍f>TMAl�l4'G�V��%f�$$[�y*¥�%X�����lw'�N�#�������kґՁ��ڑ��c�"x��n�D�%c�$�ޡ��Dp�]5���DrPE����6��r �2�.�3��	H�ZבE�z�4���ӧO�z�#"�LM���� A��t0�/LA��e`q�����w���cLT<�=w�BA#����㣢Ȼy(v��]C�7��L�4K�\'v��Vq�ὴ���p ˰�!��qwͩ�ӹ?NZ#2a��{���S��FS0��2�̬�:�2�"� ��ƺ���L�d��(_�<bH��P	�������I��<I䶮�T&�'�/^9�����=Yjֈ���a�˨Q���ce���C�m��(��V��\�r��"�j��8i�||�>�rm��˗���R��C��t�\]nT�$�>�F m�j�}F6E��!�;�~��8��[zK�Ѿ������)��#�UH����N�'Z�)eڿ�L���R�r:��h�&�1 ��������7��w�� �8��"�%5S��q��:&~�t���a���kS���������xr�u]�e�n����hi#�XUo���'�?&#Y�z=_�	r�8����H�@3USǘfl��z�p?�:e9r2�D���^7�I:����=0�u"D_��u��}Q�y��|8��:6IO�M0���nf�*"�|`Fצ�2�@d�ɩ�&�[0� :���D(A3���K��PC�qw�n�3HxNi$[fm� m*]fDH��d�LG�A�Y�,@f6�{)��%�V̰�!uB;`����V[�Q av���֖R��CNyY�^���K&Z�eK��,�͢��RĎ�RR���ȑЁꝷ�����Z/��q9�iJ)i��ꜧ�0��Q��\��A��û��ds�����Ӣm�ɉ�//˲ *�5�(M�a$
g�� ���ok�L"�M/�0��%fb�KO�-"!K�*Q|4�LĦV�%�����x���j=�m]��<���p<><�G�0璵5�-�gT=��,1ޛ8�X�nL͛�Nd��4���3�ҩ�� ���x���$��"�ʒwe�VŻx��SL�؞n�N/����3��:��l�j[�?zst a�"�$���Z�Yx�&0������;Vb�%?$w�%�����M�l�γt)
X�_�����r�[rT�v��q�%#��0`v��ط
I�a���xm�Ra�{@��N��}ʩ��'���U��y8�N�f�|��R2l��>D���:���$_�S���[�: �NnjM[��w�(9F��cH+�yh��:��	?!�]��/�s�˲�YɅ�k��&�)��	�3p�9
U��9�i�R�BRг92)%'I5��^l2n9�(B�7{��"�1�}���;>���1��{�^@�r8��ִ^.�u�F�,$Ni朅2���j=�k(�mt*�}B<��C��O��Cq㒅8X1H?a�ĤC<�7�~�B�JD���S!wޕ�9��IM�<�K>H`�g��P(��Q}mܫ7�k��[m7��CX&2QwO���kŨ@I	!���Bǁ���5�Č��"RʔR�B#�
�df�4��T��p�RZ֕�2�{_("��SP@e�&M9��4��܃I����ZSJ��D$�Q<�*@�'fr�m�2e�p��6&.9��m �o�/�qC4m y݌�������,�EL�2�>�"65w�J!
�q(X�~����x���	rƢ�:�^��7�L(Is
�J�y����$f�0K�*�ꮭB���4|������� ��^�1�ۜ�R�Nd��l|�`�+n^[mM�g�Ω��.�:�9ǬA9O�0���0z >q�C�*1ݙ��v���z�a�[�Ҕ2')�$�ZW�_�B8���9%ө�E�ӁET["U[�2�e�<=�����yN�9e���K�ǻ��Π`�"J�m�F��|�\n��5���cι��c�<3%&����b�Nޚ�˲�j��r�ꫯ����yS%�O�>��û�����׾�=�sD�GIy���F)����yRwA��HF^CE=�'4D�����dUx3WԖZ��ppH�������=# �^'�1u��'X�6�8eb&�}΅�.)�9�HT�R�&4�BB��ID�4�Qp��pr�Qy����1Ups�_���U+.6�¼�,���,��nN�u���A�0Q��2Q��(ŉ٩�!w��>���D"j����R�Վ$3mn�<�3h�|}+Z����%���Q��auA��n�wx��C;�~�����S�;s���?��'"%������M�sg��FĻ"���=)�Ku�s7�3C�^����Hə� )�T�&"�(6���㧎����?_�Cb�AA��o��X.TXRJ�tȮ���Ču榚XR��\�5���ݔ��,e�_���Y0w�$"٢b�.��ՙ*�˕����YX�zE"�/�C���-2L�r��G�:Y��
qF�c7� ^l,���GD �q��6U2��>
7�b�A���g�Kڅ�c�Xg��Yʹ�`;�\Ɣ��o?#�@7�i��,�fY�	�g�T@
�)h�"M���\r��^O��.��ښ��P��r.T�p��z��h�_�Δr�^AԃWɜ�0;��(%��R0N:
G罻ٲl"z�X�� ��"Ewg��W8�y9FWH��>>'<Q����LsJ9g���]�������������={d�Ր��p:qr��33�����{t��B�j��Ah�rA��oڛ��9�����ۚ�-�p��ֻ���DA��S�,"��SU��|[k.)��toԻ\Sm����Y�)�l�M����9�I��2y"��|8�.��4_���"b�i���ӧ��N�S��r���|8��(����)i�9	'1R2qf����Z��ͷ�~����ZURa�����)_�n�5�t�E8<]�g�I��lj��燇�)OH%��3J��M�զ�r���V�^��?���ᘧ���B�?���R�:ҵ���U"�Z1:�zɉH��sJY$���}���͝$	B��%�:G#%�Pǵ^�qwrL�
��}3y`�pq�"��B�F�3���^9��؈��P�����~J��Fx9ΕхE�9��F
��G&j��N5
,�{�����N$����|W,���M?�[�9��[�����p����n!!�C{�w�h{�"�L%g��L4���0Iڄ�z�LD��+@]��I�E8����Μ
��\$��U�6\J=��9K"�vpT\`A���M�#)fd-̌Y���e��`���e��;��9gq�H�ƛ�S(�1s�v���!�����)\�ۗ��7c��aS�	jM��X�-Vt���E����3~a=�]`<�����Z�_��̌�fZr��c����2�'y�S.󤪬���m7�Z�)c��ţ�q����+����-�
���sJ���)v6Uc!��������,�Đ��#�c}Yc<�Z�}HS5����?��f��j�z�r�Q��&�=H��ZEĪ
�Q��I{�B����y�D��!"EՈ�t�g�n1����5�'I,�LD���g�,�R���0G*H(N��us��i��Zm5$<rʜ�nz.N!�� �{�ߝ8Iw)�cq`�V�XpG��G��~����غ/v�~:8b�V��RI�"%K�%��r�Ґ;A�.I��D�SG�=�oxP��pw/c�y
�C��)C��3a��3��{oj �@���=ƨvH����~��l�Z�4��+Mf*��sqv+f$JD�J�@���6&��L[w���Fd�5L��_E�tjN�$�bBI��"��/!w������P2�A��:��4߽?���<�\��u]S�Ǉ������z~yy&����AmCL�(���\�1��%��h����ۂ��yj�i�\r�sm�6�s��̭b̨�%���k��|����C]�o�Ó`aU_׶,뺮R�u]���U�����rzx��Y�x<�pU55��-ק����LD�imU�����í�9�NF����lV�0L�.9�\��a"IǏ�d�P
E8�d�T3J�!��ŅN��5�Ȕz'rpՉ�����]�J�ψ3rH��kD;#"�i�a�>�i�
�l2�>?��ZﭟRV���f��NSb��͵��)'Bi�ȉDx>1 ]|��;�D���2rrrvmₓ�fD��c�\?��b��NaTIXc>g�Î��'<28y��ȜS.,������Z�D�(�Hx4�4+�W�1jUޘDc-�4b��&{H_���t1)l��T���J��wp�X8J/�m��SS27�^eJ��,j����y�Ʃ�w�vg��ߴ�'J��vX�D5�z>t�Gã�E#<L2m�����f�4�}����	�;���Q�X��\���W�`]{�b��P�}E��9���z��$�T�2=>>·��QO���j��@I�$	l}�M��`��/E�@�PU5f�h��d�����6��xv�V;��Y�e�)1��k�j��,*�	�`�m}A�׎Ua�JJ�f�M��H�1:Q�77rI���$#K��Ev��	�:SI��Vm�Q�!��P=�@a{��0�f]V4�kӪ}b^�;# v��4�g��?p̌�cK)3sHz�z)%�8���Kr�s%�b�<�������ɜ:~Ȯ#���jnbLf�ZY���de.d&�`IP�D�%�>3��8D����=H,�đH�)��{������)�����Wf	�.�f��q�C�� |���J�!��ML�^[#&��ԥ@@"�Ʋ�����i������Y�&�چ�f�qD|�:���������!h1��tLT'"K�H�m��J|���Q�'�v�\��ef����@��D�t�[���|��3��MӔr��HLL���ח���<?~�烪��秧ﯷ��8Ѳ,�����!�y,��)06"���z�\_____�M[k+���4#�a��(�y�R@��r7�~����x�
t��ZSI�w���>SU��jm�j#r ���ܖ�����髏,|<@2�fZ[]���z>�����r��̬u�k�U"s�4���h�A��"bI��!���3w��nn�9W�ƞ���9fq���Kz@�SӾ�aG��Z�G���h�n���2&��j~X���"U]r�9�y��|7�\$U��N�73Ws�T
؍)%��f���J ���uS��H(�X�����M��v����\R���Zɨ�`�8u ��+��H@�p$�#yd"3��<�H�Zo�5IJ���Z[�e�+��HN!,2 \����_��d�% ��:C��0p�x#�(u8�6���殭�̈́϶m�cD([>���tW��G�SUa�C�l�0F��� nŦ���-�ELwk�M�Ē��ȭ53m�֯�ZQ!
��p���0^�.ԝ
����/���qQt]������D[(��P�@6,VJ��Me��D^|H��E���$"Mۺ��ǔ������t���=�;e*��Cwb�[���//�///"����v�Q�J9vo$��DR��ȝ�ݬ-K]ץ���g�8E{�n�J��s#0bq�FX�GPZk�UI�d��̜-�u�GFt�KA8��j�ӔXRҌ��Rr.�ڈ� �����$c��ip���ƺf3�����e��U$圆b%~Pݯ�w���$IY��+�+�*21���)>��.���y̢���5RUI9��h�S�L����u"v!�C�CӀɻ$��=�Y�}�61w�4�@Ʋ�ǽ�p>3a�9�Hm@�ba��=�>���D��$B�����$"����>s�Ɍb`L� �ȅ brg�Q9�G�8u^���\�cCY����@� ۾�ջe &�QR�7��bhPɹO�w"�g�����6#�w"��8\6
���	S!�v��p�Bf|��i|�V�#�&BS���������N؏�4������,��.�����~{>��h*EkE�Dk,/3ҵ�պ\�WH��0�����tr� ���HF��4�D��Zʔsrr��B!�UF�ٜ0Z
m��(���[0�ޜ�98i.��L19����x����z���g��2��l8�^4 �#����$�t3զ,��ySM� z�^�sFS�z�-j��)Lݓ��)�º+�DbjNE2�C���=�ugH\�uE9�)9�yr����!"��ڥȼK�1�sQwkJ0Z��̪���({+#�4s50�`aa�oV���U$��kX�ѕ"�)	扇���w�m����s­��F��}�)
 ԝ.E��N�p��m���0��)%I%gU��)�=0��E(	�Φ���+�/u���LP��؇��E�ox�V+3wx�U�����^�&��p�
|��&#�9�Z�ӻ���$m�ܭ��Zkmk�	ֹ�2;�>�0�$��g�|q����w[b �����5�0�X[P�6ŉ`?�Gg�9]�,�<%$��k��Џ�����$�Y��x<<<����������v�9��<f&&�&(�p˲���o��W��烈,˭��Kg{�͹���"���벬�� �B=kq'�L�=X����df#�H�{��.����u]S���#HC�2N�tv{�M&@"��Ak1w���k戼{_Qm��VH�K�_��	�@v��8�5������ֵ6<0٬3(�B�e��p]VGn�K[�"A!&m�cO�v��:�%rI��e���u �Q�R��B�h 4hʡ3Lv�pS>"��֏�+�c ��������Sjk)oX?��)�\��4��@	a��=%��s�互�d�,9'��A�]��8a��GI�EDR��v"��� ���F!�����%�xo�a0����x?"9t|�+��։�W�g����#�e�l�y�y�R�3����>fv�^�6fι��}m+'��̭��c�{/�늽���u]��3v��t:��d��c�f��,���eY�9�Rvb7��z>�!6�}�+ǫ֊ɺ�V"d�(|u+���m�s�MD�#�r�}��9�P���0jq��98��C�T-��rk�"�-SkFl�T�y*�pJj�Z[�z�\B&�Q�4���̬��!�J%�i��|Y��PBEO!�eM[��uuT�Gd-,8Q5��c8S=L���m#`"��b�hcωo3���U� ��AS����{�S��*�g�	����'�
��&����Z[�������3�n��HJQ�S�Dw3l��F�;��ѕ�W��
Q� -�G���gPX��>����"D���0D�Y��݈���uiJ�"$���O�$�Č���B́ݠ&���c=��A�g��nSE��LI��ScC�?��p�< ���B:����(�`38;�N�����Y
#w g�^�t��ӌ�f1 A*u'�!�y��#77��R�D����yq!cD�����������.�tlw���.3w3���\�4թ�i�J)T���!z�] �:P�r�u�y�?|�x��ί���%xBB��͛63k���<�������jm���p�~Wk$F�Jծ���z^���u�����hs���IR�3��R�K)9'�V�Z@
�hM����Ţ����mϠ�l�RҀ�1�Ωik�r�0S���"���j2�4%%j�UwO�v�����k5�>>h�[ ��!w����
�Ȗ(*9��@�W���cϾ�c�)m�3LA�Ɇ#����K�����e���?��A�����.�ʠ�	;)�NzC7
�{I��TN=Wq2g��XR�}����J�h�����Nf�?{�f
�O#�U ��j��

c/H�{�����ad�hvV@��Y}���F|��ܭ��GM�@ID�̵-��q�;�~p�k���X~ۄ9u�X�P����I)��������)N=�*6���5E��0�t������V�k]C!�����^>v����R ��9>6�6m��j���z��Z7U`3#�RJN	 <j?(�Ѻ��zSm��"��:F��������$3��kS&���u2o��0������L9;�	V�\Zk�~8��<��g]�秧�^��e��q�GW���ົ�}IN�K&����S��Ѻ�]�f��jj^�5K��;`��K1��;	��7w����k��<9��nV�����[�=��Ok֤AA&J!N�@��Q2����Ff�RFT 6��"hF$�����E(,�@&p�Z�sI�����QҾ��$�Tq�;�����=%<���7��y��S�N��I�oQĳ�8(:�$�Ȉ��)����l5�X�s�]A����n;1Nx��w�2�e�a�����Ϫ�S��[;�Ax�镰9�c��Bu�c�f�f΄�^@	�+Zz �B�FIB����D�Ams�9�0��#�"�M<��$��?���U"�FEaA��߹QJI���������4���St�pk�U[��4�l�]��b��P����Ø�nK��x8><<,��֚K&�u]MU�����07�������t"��ֱ[6����H*wr��<??��<׶��K��|�sJ� ,�[B�%�C,N_)���D!�Ć'���\`p�m`ʽ�a�E�Gr���Ci�Jܵl{����ý���P�׽RJ벊pJ�`��������=����e.2�X��Hw#�-�5�0z't<,|Qk��,Iڪn*I$:6⌉H�$,I�Gy���N�\1~��M�7��w0�����BQqS#"'s�c���D�������72����-h���Mv615k��)h�#�vS"�^K43b�����n?�pw!wr�f���X�
�/�v[WSL�A#�r���ٴqc!���w좞n9����h�2��u����P�#壆~��E��ZS\��u+Jf*��OoZ[��Aĉ�i�u��嶬��<M9��m��3�����Lj��o�6v���OO����݇i����W1�����	t#DlI~|�$ɥ�6�L�� fK�������	X!�\J)ECa!�QIE8�L訫�1l*Q�BX0&�<�ʔRau_������|�k5�R���n��6�YYN��nu��l�ɚݢ,)�tY�RKOֽ�¾Sw`-L$ν[7���M��Ю���n�q��03��I�q��0Z��� W@��u8T��1��������0��N�/S"��� f*��ɬ��V��Zc�*)���9h��)IJ;p;���������SJ ;�uy���)VK9,8�S�>c��������X�NL;��8
׭E	#�G>��pfiM�=g�>\;��ᑛ�z0�wz��1c���E�>�co�Jzw��Q�#C�~cD�����(P6@/Ȭܓ��D:�N�A�u������UV9��Z�Ʒis�.�Y�q/Q�3%�i�>|x���{�9�Vk�^/��e]��sOބ�['�"��);s1[2����N���2�Wչ={w���r�͇y������r��;�K��,z��i:OS)��u]���Y��M+c�@*�$'m������r��	d�A�6D(�ic`�RN��4M��6f.9K���z;_����Q\�N��s��z$��8����خA!�;&�IԶ�W37���3���L���u��͙���ą4��j�Q��.��鏰��(��L�ڴ���Clww���ڰ<(�8ui$�`Tԥ���*�A�y`�K��Jׇ߸1� AEv�nn^��D�kn�l)��D�A�N@���I�`{������E����F��S��]����m:��0\���!�����hK��	�<���Сw7S�v$c+�2Ww�#��]����z�����@[��	���R�R�sPS���ܵ���ߣ!@MED����	��4f7o�����p��yY����Y�^F?nl�G"�a
g��Ջ�/���u�S�E��S�E$����Z{�'�,)�����֚����E�q�ߟ"����_r�j��I$��QXZ���3%��e!b2��J�S�,�w�V ۰GfƐ�'N)y�y��ݫEo��ܾz�����M��w�y����&#���ɜ�i[�5'�x��C���ОƉ�t:v:��p3�P�B#��>-R��^!��=�ޟ�8~D$�:�F#I2���:��w8�鰿�"A� !�$8�kn?\-x=B����w�a���_½��=��W�a3��������`��/J�����֪��]����_3�3t-��G�|sa�1�p�2�I )z�zH7�ߝb�n�)���Ջ���]��3_B����6
�=a��fǻ�;w�:��ݫ3n��R+gՠ�wEw69���� ���̭Y�MM�%�k�����x��#*��v��˷��% fu���0Ǉ�w��˲<==ݮK�mYW𖰉#!F��1���c�ISIErɅD\�j��}�9b�~��H���l�*b�ٝ��x<O���޴��s)�y1KN�r.%c�vJ�,f��ö��IMk�)I)�����z��/����e]qi d��EJ��D�����Z���y�&���$i����v���E��G�f��A���?�~~-(!j�_+w�e�$�T׵5�'�g7'�1��I0����N���oѭ���n�r��ֲCz�R3k�\[M�?ۙ㈱�Y���!u;@D��6m�_���s4��ZG�*�5�wn	��	�@���܌�\��̽}"��	�Oc��ҏ?��n�:`�6BC\J�>�!s
q�q�}�%��d���b_�%�����Z��!<T��>a��6f#0Ehݿ`?��A�9���f���m�H�&q5��i�m���
r1IJ�y�4~ a���M �@h�~��7�뵔r8޽{���~��r[Ηs]k��Dk]}]sN9��QNdAVo����"�V�Kb1{yyM)?<>�*�� wRl�l �����+$+kU� w��g��\�eY�jfYQ܊�E����$�Y�P`&¦�A.�H� kԎ$	H�fD�#�6 0�,"��r>��7��""���H��As�����7���'
l���:��̼�v��חs"L	gX2s�u���E̈́�c!���;y��3��(KF<A��¿��1�{HG(g0� �oh�ޝ�S�)�������cf�%:�g�m��p%ь$��ةcZG�`P�p��x�������6x�}��D%aւ9$���2��fNĄ
�����s.��"{S���#��� �c�X�F޹/�Ǩ	��q<Ia��{���~��l�>�����̕���\G��W	Mʠ�%.��J�Tl���:*Pa
�{�Tl�q��D��_z���4f�\^o�k���?�����z9��_�|]W@@�����䨴�Ыc��97#5��s.�d"���s������I�,%�b
F��eEK��p��m0�N;9�$e�N�S��4M�"G�؀]�{�R�T`�ٺ,�����r]��#��o��� s#�&�֚�T�ї��R
� Nw��rk����;w(�g �؝�γ�O�3滰�ȉ��;?�6Z��8g01l�� ��)��o�j�#���4R���pgS��ff��Z�CoE�����/�Lvw�!��S����2��x��q�����(=̋*&<z����JMwLZf��)����A1 wO�E�?0�q�73g���
��̕#�·��r�ك�&�N��XXH�������!d[�b2@�+Q3�{(X@u`����0쯥R�͆���G�ΉФfko�����0ʡ'x�9�����G2#VK�Ҕp,_^_Zk>|��TJyy~Y׵ju*�s�5���j2�3�>�9�	�
Ѻ��۵L�4M�*�S)�-�)�;�Q3ef�4��-��R&Wo�
��+w3��֜�T[�I�Y ��VJɴCȼcYX���2�����D��̼'PN�h")h�h.�qA� ��V�_����Q~�Q� "��T�t���;Е<�d"��j��Sy��=���Ȑ�G=~���9��䣈�)q��G�8>��	;����C�E��.�#���{�*����~�KG�8x�=��E^+[�`�JS	I�N���G��@sU�e�8�Wd�@�WݒҰ�Q��Hu#���%rf�Q�F�@��;H!�	����ْ��"��S�
z�to�Bjd���F��n�*`� �̵7����q'#�ا���h/G����c��:D9��֤݇��{�履������;7����9?ƪ%���:�� ����"KwN�w�\7�,�2��,˭]�p�k]___����1sJ�['Ǹ`3DB>��ȭ$�i]sΧ���U;�	�?��j��8V�!�Wk���R����9R8u����q'�@ѵ���4�Ӊz5s]�����弮K'c�� �ys@P�H�J*I�n�r�ި���z�E�c	3���H�^;���I*D(����7ܜ�����"�в�P�uؔX5M�9�":�g[�݇h���t��HȦ\���]'�\Rd�f���|q�1��-����R�{��-b�;VE�Cj.~�Q��e���0_,�I���q$�,�-ر�"A��Mɓ1R�Ѳ?	9%��P�[��J�p�)�8�Ѩ���i�O��ѓ�bP0N���29��=ְ�/�93a���Gĩ��{oܝ��p@7$"�����/��x���_"�\
��p�S',_����#���m]��|�_�e��>��V!q_c�.� ��zE�*wU/&�U�%K̒R*�����
�g�-�r[��*��OS��N�p�x��F{�C6��v3�fa2
���	���:��f���l�F�ܟ<d���S2o��b�A�����Wk��S��B@�#9�U�e������j�)��=�Z�L[c�,Af;������B�TM�e	���u�H���Ǝ��.��hX���آ��X��=z 1Ḡr*���R� <R6@��c�#�$�n���:Y���Sb��e�1d�'���8�"̷�����.�$�N�W�h����A�d%>���h��nd��ǡ��_"�	7�cƒR����T���}��$��9%�_��l���LՌ��xJ2��5C�r�齷,�\Od�N�mBԵ�;�oC���6.��Ƿ�����^܉��[^ �orN�D}Awu�0a(9����0���,wV{<5��.Bv"��W���h�4�����:�dC�m���aQ��9�l�d܅��v��UD�b��f��Br�ɜq�RJ��4X�)�i�p�q���"�uYǟ���r��U�y��|���c*��"��\.OOO�r�{��|�'��2������<'�IyL����ff��e�N��ݥ�>}��o!����cڍ��$N��=�EH8I����l�h7�}��B�(e���Q��&2q�JDTR6־s`�d�naJ$��Ș"���7[�,"#�r7SN�ȝҐNE�����S���: ������S���v�]?��N�7��i�S>��-�o���F�OD�6+���l΢�z�+ ������ay�#�t�εa��8�Yyx����&�^�a��w���&��h�fa�SY�{�sO�'|UO��=��q���Ǳ���g��|+<J�M_����9�j�n0�c�!��D]W/Y������)�|]��9�<��.s�Y��Z��A4��y�	"2&e�7"�)s��O��	�ip���8���{<{""�(6��M]ۋYr�s��O}ㅿD��],�Z��&q3�Hs]����˺�?� �&��M��(�����G���'�N
o��Gl�0�u���6p1~n������c)��=���r�h
�#�[p'J�b�q�f��p�kw(��ɐ�d"W��$���려Q��/�)FW���N�(E��[(w�ah�'ǩ�{��+iƛR����(�dcG|��p�m��灸Ek<�$�O!&����,L ���0�A��	13��Ƚ5�V19s�O}ڵ8l�m���������4m�U����� n
��&��.��.�>��������@��v��w�2ݷfa(��\��xc��Y�RJiY�����뺖Rv[�?7��w��Y�OXƩ�Z����u]��<�8����w��b�u6�}tܰ#��N�%Oer�T�z2��wuI)s�55ss�.����z���R�2ە����=,���s�m"�ۏ�L���' �{����3�㼌���h���㡝Y���NV�6��,������m�?J�I� �m���a�I�W�O�D`��K���u;ܸMI��:>	s)���m��g��ڶ!���K��́Dz�nUH�E��O��n�a���qw��_xk�=}Ӣ��W`�ob��02���x7�o�ܻK�HX�+��&P_�q�9�� �o!H��{NN�/?������$�#���6�D�������l1e�*F��D���6��+�� ��Zk_�0�x�͉�ڲ[����^�8���z�8UsgWW��jJ2�R����	}�{�{�]�����
��j�=rw��R)�r�	'wʒ3���L���q���ndj�ڢ'�w55�nծO�Nn�x����P�� ;k�}G�5�6tVi�߹�u�<a�y7a4���C#�&�7"M_��%��pꙚ���Vڝ���8�� I� =�4 U��rߜ�H�j�E=aDD��a��>�`�H1�[�:��=5��������+�ґ����m���{�ڇsٯ+×R$�#F�_����2ћ�`�)KO����P�u�]HJ*�d�L܅��`�np�:�����۷��H��L9v`'����Bo>�9��Q���)�x�vf�h��h����-�.g�[աl���A�vg�i8N�=�Ǒ��kУK�Iu��@}}uwt}"-ѝ����m��(c]뼈�%̌��Z[K�:������l�&]�P��1�����,V��.aX�W�0�yQ43��L�ֵ^�����%kT3Fp�x�{�x�}�M�����QG���e3�����敇܌�>��u�m��g/���õ�οÍ�v���]t���h_��;tX�t��tr�+)����9�����Jsf�)gw2t�n�����8�8~��	�J'���� {�d��·n�G�Eچz�	�,8�w6��RX����[����f6��%% U	�x�����Q�ض
p-wB!���n#�}i6'�_�=�M��>������������j<�ݿ���U���(���9��$<r	X���C:6�$��}J��)��P̬���D<co��;�"�mY^^^N�SJ)3C�=�K�.�$
r�����Ț� [Dzr���#�NBa!�M��$���a:(��'�}��!��������7�mؒx4���n�[m�S+޸<�38�����_�ܟ�� ����hfd��o�h��˿��Ѹ�&���b�D���z��tA��n&�H �<�ݯ���/���a �l3�9N�Β�8Q�c����?{��#��R�������(�7mNo�bC���7��>6��O������{o���Qf�!�G�0���_W�y�N��}�߆G�{ؠ�'$D�AІ��$!'H�w��LԂ�Ӄ��RlSX:U��_c?�!0�c\θڭ?�	d"D{��1��G�qwF��=��>~ۓ.���DJ=��Է��i�
@�"���q[��T����k�'63��=-'"IФU͛ݮ7��\�DƘ�q�]D�k]i���Ms�US�خnޚ^/�����*w�C�����A�t��.���e�L�35Uv��H��'�p"6u�Fd"��}+�.��uo*}�H��t�AC2�;�f��쑙�����>����<I`W������8O48{�1�c��l}����%,*��T72��7�����������J1L�o��$�駌G�>��.�£`�R'	c�v�Q�7�{B
� �+5�}p�;c#%I�4T+v��B!f�)c0,���=.�)^n:�7�k�Ͼ9r~��C�)3wFmܯ۰�]�)�4��;�q/�^�hcr X�J�����*��3�v��,�/��p�b�z$��b���]
����bL�Qs� ���H]Rr3mz>�SJ����A,����ɛ["N,k�[m����UBL4����#���)����JJ*E�aP!�Ti�JĹL̮��y` kN��ND*6�%��4_��T���ٺ,�5���-w'n:��nyeۍ<ܻ�$w;��8�R�m�Ʌ�#m�bV���S�����6�Po?�=�4�I���vh�;!E����1�X�u�V2K0��;9�Z��]�n�h�]q���~qw�Cc�G�������̽m���w�&�ʫ吝[�o���`�Dڒ_����E⛹B͈��B}'J�Y��U��nU�n7�Û9eز��-c��BJDd�vM�0p��B"Bu����z�mF y��7iý6dWRJ��$��4�MW�=��6�<�3횮xd(1�b(��7�y�*�]^!}���69Q����즭���Z��(��j��2K�)��=�-�\��p�F��-u�2I�.��唑�E8�B��<K��j������=j����;fwv5���ՂO�c�,��MWEK@ι�T��Kʻ:�>1N L�Iú�hf�͢l���1NΠZ	}��Wą����{�w�%��,ow��~�� ���D�֓�}�	����6�s����.��Y��Q_X�����.!"}x��o^�AY�þxØl��"�[��|��-7�-�އ�� �ȝL= Q<��kL(ۅ�:�����n��;o!����0w�<l������ �Q�F�)圓6�|@x��_Z:=�[�� �Kt�z��[�曕��w\�C?��Ɨ_�9����IS�D��P�";a�6���벴Z��!�z�imC|�C�s�Ģ�F+"���X��I����nI9��1J�MX ߚef&qr���cxA��B��خ��P׌�SN�CJĉ�6�16�[�y�q�-�4���C�#bΞ�y<H��>+��qa��DtVrG����"�q#��ۺ{R"�FL]
.�����$�`6_;.5�f8"���=��8G<P�X��S�_����K��W������������{�A�����V����ٌ�v��N��}������EVH��j����![��*2љ����{���ˋ��7f�9$�m�`!��?l������폰r�������=�����%��%FC~�j� ��{p��n3�c4��a�"=�N�(��m�%R�-�!~�ct�jӵ�Uk�"ѡ?��Xtf�\r�R[զ�ZK�@:G��{Ͼ����l]+A��"���5զ:�hyt��L������H;����%燇�e����v[�[k
���E""���	��)�Ƀ�����0��-����٬I��ػ(���o��ݬ��'�<����en���p)_x3G�RjMMUDxz�6%�'���"����l�|~��wwuG	�?S��d�D[O[��� rwT����'0��-��k�F'�LAg�k��Ӑ*��g��㣻��r\�y��;�>�t�ّոS�
<3�9�]�=?��0sm���lL��'��m�2S���17�YRB�@�i�f{9�ܛ6b/93�Bw,�8&��'��kN\��63Ń�^�f�^XXU!�D.�.YDs"��m��)cUu��<64�?}'	�K=�!��4�Z]� �av����<�a���[3w��K���r�H�{���)9�u���c)Wu"�D$�ZФ��8F�(�;�	w������/��������aREd*���3wO)ńV�p`̜���#�n���I~�p�?�bB��Lͽ���=������{�f�������(Z��-%��K�c~�ջ׾�v��������3���>���y�"����M��/-�4��v�)��w�>��y��<nb�K�Ի��0�����ݛ�D��B�)����\_X�7��Ѷ�wA��owh�$����S_�=v�w+t�ۍ ����&Ձ%���`�Γ�?�n���1sb��S����q`�9�$����N&��N���=�&��,�q����[f���W��t�cΓc�EM'�����R�i^�u]�y���n73�)C�,q"�u]�Z)e7�9���7Sɹ̓�Y5��pk���@\AK5o�643�����;��?|�p�����ۿ���xzz�^�����p|xx�9����v[ֺ�r�8j�����/�� �3vv�$q�v��w�{�?r`���R��-�i�uD�?���}���i~�k�1Ԟ)�B��=N�8*`!+d���u23����nK��^w�-��F[$���9��o�sF���@�"�����#�l�I�6��.���92�7	�n��?踧~���GcX��MP���?c""�;�e��v�jojC�t�p�N0!G���D+h���n�#��/����̜:���(��?�|�r7E�hJ��j�E8���fF �fJI{Y�G"���@�9G�2@��&e�Fh}� �5E �qS(E�@����zk�.n�S� 4���7�h��.3��36|��Y�ۈM����O4&w'g��w�q�����[�'t�¾E݉7 �P��~��w��%�p��>S�S�a�saQUf���hL�����+1puv���Eh�f��f�{�����F�Z1xv�~9[��G�\��c�-�G�W	��Ϸtd�P�y ��������+%6gV6��s�~7[O��JRD�a��M�z���?�˯/ܬ�����Կu��6��^��+���vC0��ـ�p7h.���@ۙ���jTí�|0<�b����0#28\ޝ��o�OB�8��,Nc聧2�?'K&�-�Q}᮸ԏ��m��urh��?���)������|�m��ٛ��؀I9qcS�Z��2�)Gj�y��	ƚ������3M%�<���z���a�zh4���u]�՝>��x�O��痗Wf�T?�Bj~:�����������������_�����~��L��IM��Vtq��N3�d&�Ҝi3Sb��ɶ03��B�]K�O�!m�<����� �s!ޏO�â]T����{|���7�o���"����9'H0�E:�N`>���D���"�{Ǘ�J�c�1]ؔ�;D�M �}��/����x��-&sڑ+�͞W�׶�!�Ɂ�t������v(�x�����w|�?�7�}w'��tW��0Cpi?-e��x�6h�D�D�; 6�'\)(mo}��� ��{�B#��s�Gd f_^	�5�Z�b�MȄ;���%a"o�Y[��߾Y4"�rLJ��� �R?~p��������M�P�q�ssr΍8��HF���B�[��U�w7wq�����D�A��K����m�N1����P�Ϯ�_�Eo7���g��{���}S�'SN@];Bx"�%1���j��+��>�S�E���h9<s�C|�!�"�f
��$�C�pǠR�Sta��D��tk��ٍ��1��]0e-m�2���ԍވE�<���ya/���|��u�!��#b��>�f��nw!��㟇��;���]���p��el�����w,��Y/�]�w|��A�o���ov�$L/Q�c
ݸ/<�/�h|���	�ݻ�_�����Tu#��b������E�w�9'I�#��ޔn�=��E��ag���ѣ�E��5m����������aSkk[n��x�)W�j*,�C��4�r��a�,���	�o12s�7�B8���{8������o����v<K)ȟ��@�-��)������������O�>�iBA|���|X���JDY��W���M��iÍ��M'�t��D1�·��cF�%��4�Ę�Ń�E���ZC[tkcj���2k�#%�.�;���P�)v&oJL`͊`�����|4����j� ���S��^�]�Qy�?��
[��sgI�=�L���[�m�`G��F�96�����}e��7@L���������C�E��h��sĖ]�?�����lw'G; /��΀3u�O���f��3�-1����5��A<���w�r�j��7$���š�2����Q,��J�#�ܔ�(�g݊�kӑX��6�$�����s6�|Oy�,1�X�Ӗ�'e��E�RJi�w��Z7�N���]��cY��2~�DJ�lL�YRι�4���0Y�)��%ܝ����/۸��%,1�7m2�#S�C�&������J�T��y���y��;)~\ Q�����,�3DD�䔉xmFd0^�)tGUU[K����E�w޸`|��b�)n*���f��9JcfL���ZPSbf�WZSL
Dǃr���J R�D��1��'�Gͬ5���LDͶ��1��� #�A��o�:��<���r;�(��I�D���F̸?���_���aP;�-�Wr6��O�;���ط���Aw������z�ax�!��ştĝ���m��-	������kx��K)̰�u���q��������O�͞oO�zB�!փ�!��:�j�}�`� UN<��X��_ R���_�y���is3��~�_j��(Φ0uq������q�3sɥRm�]��Rr)EMU���i���BD�j�f��Hj���i�=50��Lܿ�2� ����3���'/�M��|~������������?��O�~���������)ɔ׵2sɳߩ;�ϓ&'gWS��l�]��IX�NȦ�&�o��v�w�ߐ�g���)�W�hUu�&��
f�$	�)(%�Ϣ�=&hI��ʹӵ��Yk�1��p��W?H9���b�1Kk֗��J�$	�1���^�Q���i1�	́@Y�<��T�YߑF����~��#�o�{ř����!<E�!��x�Ⅳ}�r�m|dAF�E�������"�!��`	ڠ���XB���=t��[t1VcX0[׶5�d&I�Ǖ���Zm����� �@tm!�P} �4�$80iH�q�ٽ-ˍYr.Dޚuڷ@���3�)��ڪ��i�Dph�Q�q2�.G2kx��Ŗ#�ν��$�q���	�s�_p ��}_X[�<�^$�OtGΎ�)�r��_�lUD��(K
�n�^�y�����=q!���XI����L!e�-ƇÍ��a8�h�J)��;�C�MD>}����;@�벮����T �����Z���<OLn�Bb �e ���V3O�)�ټ�C��i��#�q1&u7� �y�rB
efIR�"v�����Ġ�Ũ���D��SxUD�)eaV���#
ӑ�D���0@k�YX\t<�sI3�)��;$f�Y|��D{���Q��},=
q2��Jê��RNhdI);a(_�G���c;c�d4ZT��n�ɸ��eq"�m
�3��2��[ll��nIY$a�wZ:3)�	�;�ztEؐ���|ğq\�nD�j���>0g����73o��FQ|�e�a�e�"n����3�G�Q��l�w75�H`<�ld�ֱ��[�y�Fǟo��! 3�P�q�"w��C��)I2bU��E�S�`v�B�G,��n��ֺ�z<�LM���`ڬ;�m{���s\U�)ά�ΰ��`J���9��z[!s��~����|�uu'U�����s7b��$��|������������������?�����￾^o�D�f�	l�:jW�M�+�M�93K���2F�y`�c�zW��	���ɝ�SH�$I𢜘̌C��2�4#<l�D�p�8˺�p0fА��H�Iʹ�\�G�j��������dd�$f����&R"6��.D�<��͚Hb��!:'���%���fʎ�:֙�̶C�h�!sW�1��> �+��Y#�2�:������w�9>2Xff�j�H�¾%Iy�7�H�ݭg�q]8�þuiUA�Ϩ���c���X�{A�a�I�S��DIS(G���.�L=�Tu'sE�@���5�6Bլ*h=#j�}����ښ����Pv�P� '2��*T;a�M��9�5ߍ��E�ԍ9����ifxվ��?9I$��Ƀ�g�dd*�LfSWաAü�(�=�aW5� ���$���a"%%�ഺG� ��RFOja��A���Шs�sDD��������k��&b�����)�]攛����������>�NĤM׺��J;VK>�Tۺ����>���׋��Ӳ���R��u][����v]R�)����$FH�K��-���<faq����D)f���6������Vkm9�X"��,��|�2S?!ԕ�"RAc
�PU$�UFa�+��63�3���Zk��M���Bz�;�а6f���cۻ�9Z\q����Dh��!��Z�r��%i�������|��No Q��-�~-��G�X���=�����45Bt��&I������VE8����u]F���ǫLSJIv�����*@ aO)#� &����޷�D,�D��Ͻ�),M��!���@��0|��L�-ۃ�Q@��e�^�����y����=j։t]op�5ai�p�IpG����J�)e3k�
2�ZmZۺ�������K���^�1ȱ��"* ���l2���c`���@�w��Q�:I2�ID�9��,<MŹD0��`��9!x!�����jD�l%O�á�*A[��t��d9~��_���O�Ϳ�7�g����	�Z�]��wkm�m1�RrJIuE��s�織	����U23�l�,�0E��c��H*�C�ϰ�M8�J��+2��KNB�j�K	� �Ӕ��8���Z���m(�83��Q%����s������w���L>�Nn����.�<�Rj]M�LSN�EB*%%'J�M�HH��%"$�AGqU3M9'�i�}��po1�1����[G�����8��r��o��ɽ��E��P�P5	�~����ͥ��+WUf.)�鉈HRk`��vJ�I:�Yܥ�;�j�e�)�aN��NA��|��x���H�ǭ�ր�&4ћ�z���S�9�{��	�����
���D��ΒJ)�i̔r����w ��$I��;�pm��KN,t�][k9��2��f�̩��n�u��T��\kw];��F��!vB�7K���?���r��5S�>U��9u�����<�O�- ׉g�"��U�jӖB"Y���qe��+S�1ͤ�ق��SI[:��B:���119� T�]���w2�����2���?�я~t>���_��h/`am�֊:�>~��Tk���~������֮�����_���q3�TE �Z4�������Z���N����I�1{�j��J��km�mu��K�I�jS�$,�i��!72��`��,�1bq7�N�Ě:���r.9�p����Cc4VO~�Y���4��ua�T!b�Z[�mp"b��T�vn���o���A�|mX@��}H�G;��$���(�1m& ��?B�ɕ�%%�Hܘ����p3�Rt|�(W)S�	�UkU���X��ɄL	c���AK�r��__k[U�]���
c7Mӻ���=>�P�I)�R��L^kE؇Z�%I��ZW7�$��Oh Nj�c<�	`F"�M�6��p\D��z�=j�A��2G�h檊�����R�,�]9Kr���� ��W�6�=٠]��	~gG�-	���t�-NTrI�m�-OOO��gr3W�"c5�e�/N�$Q&m
ۺ,�<��<1#MRi)9h�;7�۰��qf��������ȉ�ik���J�j���M��N'"Z����i"�Z+rT3��JDe���31�n+���pH)=�<������N)�ZSu�̄�N����n7"��9��Lj�b��(S��I�� �s�aK�J0�s�G�HO �u���8�,��q*%� n4�u��~8�Ld��<�211��R�nZ׊N��.˲��Jg%Ű�V6����H!������?}Z��朦y�`��Vk.��4�Z�Չā�D>D-�s)�$��{V,�S� {�E#���,*K�xq�b[�p
$3 3�9�n8�D0�¢Q�'�'yXB����S3 @�)�{�5Kr��Z������*��4G�PMȧ�9���ִ��2Q��J�Sp��޳�[�.x	�@bɹ���{$�2Me��	A����<�Z�!>��bށ�Z�#��`�k]�HXZ[Z�eY�ur��t]W�9M�t8�y�����Z�P�d�GN�.Kk�mӐK&����Z��y>�f�H�i]����W�W���_��*�q+��x8�p�n8w,�nb�S4K�G~����V��T��[.�3;5o[���x\+bX �G
���%kT����,�Vf�(.&S8�d)}p�� �������9��چ�R������x���幰��m��<�(�	�3���c�n���p���<<<������o.�+R�$�8������o�VΩ������~�U]׵./Oϵ֯��������xć�Y)�p8Ժ�Z�3/�;q�j6���|[��a>L��wߍ�q_R&�<efIs�s��,���<��~�9���u1�fJ<&����"V�#�?t%��{0&˙�(H�ú�C��Q�dbɉ�A�TQЦfw33 �spw&P�J"")Z��l����Q��ZL�.A�7�O� ��i@�<s�)�Ć�$v���r8uf|e�ٚwzz$d}\���y΅%�[ʉ�km���sd�N�� f/��Z;��"Қ�� VYh_65����n�=����{���������@x�R������Q�k5MSJ��.���%5�4i Ǒ<���?�eĩ�?A�U�RθfN����N�����rʥL"�)X�]3^�ѴDIR�$$(#�G�Om*��@�Ir�>}������r9_����.!���ވ5���$�kmu��44��`�Tr.h1�n��x*�/��ͅ���\JQ7f/�p<���۲�j����n����̏��Nt�\������^__��t:NӴ,�}�������)����'R{z~������g���믿y~~)�����%�q]�4O?�ɏ�����R���}��7?��o��'?1ӧ��������3NI�����8�f�)��S��L����I�8*�l�n�������uJ�9�� ֺN�4�smU���R�`X��[���JD���x<hk��b4���LL���k]k\���p8�<�����z1��'�t:=���vk�F]GP�L(J �<1Uk���|P%�G�s����$�X�3I�����m�Pq��9��CB$*w�����v4�Y��Ro�	�09D��c��I�p9�@~ML�j�K��Z�Z��ג����ZmfanW#��&730Y���{�SI9疒f��3�k�9�|9�a'U7�I3�ʤ�/�/�����y��e�F��|^�������ckM[�\��Y� 7���̦iz|��R�7�֊&x�)璓�����4�w8[o�C)UJ��"(Z�ޫ��F���[�=��F�Z[��B�j�(j���V{�����r�:����}��~Nr��T�b!��� ���!u�L�=)�eg�K7���w8Z�/|���d�w�����x	��R%���̄� ��̿��)z�Vf�=8a:��E�_T�I%�������{��D\�5����s�C���^�!jk^�y*	����Z{̣Fs�w[�]t��	�M�F��K%P|z�-cyv�Z�>LH���E���{q���{"K@������ͦnD~OU�>m��~����A�ib>S0�mEі~:r��ߣ�����E�(w�kj|o�a���d��Њ-�1��Q��8*���f&���F�?"'/�	:\˱�w��1ljoz�t_Z�~E.ſ���JPh��rV�>�MöT?�Wed$$����� ��š~����h2�-e5��ז��q����CJ�L�i!:Y��q?js-:�d��0#���������S𣣢���g����u=F�_cw�.�nѓ˖Q��XG��>fv���2[=Dsʔ�˛׶�i��ץ�%�
V�}?�)�Ǯ��������Ҹ�8�zfo��(UO:���^%�g^�+>��|�<p�ro �٭"�G���������  �t�,aq�&�N�4���)V�3�/��h�'���I�ԹC��(�����ʕ�]���93���%Z����;a3�a�����`d���bGDJ�Ug������XL�왹h�b��h�WӋ�_b��eq�+%��[܀�!�=�+!<Nj��ْ��PMB3xK�dZ��/�A���J`Z5�]7���n!��m�X��yuF�]�<�[�^:MNa�^ ���rW�]���k��ZZ�o�+4���qPs���'��5��t��"s%5��f���9����	Ѱ�L~��i}â2�h
�5�I�Bd�oNN�R�A_+'Gء��Dߢ�%]�Ni�� A��b�"P��u��c�uuf��,g�����sU��~:��XgL�[���KK̝5�|�'�ۿvv���������z�lBMe��v�UK���V�Sf�[/}"$�E���7!�� ���>��esm���adF�&�# P;ܺ7g���1�v.�M�h�l4{Y��U��^��c ��]Ko�S�����i3���o&�(_�Ȩ�BQa!�|��hƐ�'2K�Y�)�)�i+�r���!�^�u6��#�����,T6	���gT�o�XT��#="i����Y����.2�M��OD�d�O�b��_-�;�.E0�{�ɀl?ƺ��"oiGſ�+=����,RJ	k�1�f���J^���T �bڛ�h:��b1�}83>�a����
^b�����A�g�'T)��g�?˅�BvY���e�q�ך\Q���t�X�l�^�#�ק2���Vim�dfaYl��[����������W���Ԏ\����~����b���Ѯ�ȱ�<���.��\^@�-���?n��Ho�-K�P�,(O-��9D����J�Ȼ����S|$N��i��GO\Iu��q~�(���O�ᆡB��X�H��C�,h>���$�"�w?��L���8C������3`��O����=�zkn:x��l`�X+`��1��)���98hz�O�NS��! 4�t�Ke���%r�F�S��E�%EP?Q��DC�ɼk���+����=���l'�ߒ�%0�u砲�A���q��.<�����������Q�����LK��|�Y�V���E �J,���_����l+�)@$�Q���[��7��$�#�d=�{ll���t0����UZ�����8��Q����=-=��D��l��?���҅���@����Ն5�<�������6�7��jLN��{���O���YFکƨ)���҄���6!^-Q=�}v�_3�Fb�W�,�}�.
㹤�G.�7���[��0��%�hc���|��	�Q��.���!_�Sᦴ?���5�:sǱ�6��6Q������0O�"Vֈۋ?������(_ڃ��o׼�6x��lB���>U��p#|�7_0u�� �I�p���v&�n����^��>��m���@�؋^��2u�����?x���J2w���|q��������<y�)I�6?1�A�3�8�K0;<p�fQ>��ޣ�7�e�Q�\��[x�ڻ�P�s�`�r�`l�=�����zB^M-{�5�<0H/!�����r0��#��~t��j4@g�'�ٯ�J` �F���F 
��ё5}��]���2����6�������~*e�NnoLp�~���M�U�������)n.�﮸�J�t���֕��{}�����3��j�/����#`���xI�u�u赗�P���ř�`���pD��g�/���A�t�T���hq��?�6�����w�wi(*�|�� ���`��Z6��8���`v��#2Rzj������x���3c?K�����vQ����=z�",R2n-�=�x��z�4�*p�͙��8���I��w�����H#sQaq%x``�x1~���l:6#cř�I7Y�_�o���*xZ�B��9J�k6�S��i�Q�ѧë��:�M�8�˯z��!G:��/�`���#WrR3�����D�k@|��!��)4?���^�J�NH����O$����G��.$���%����`��C���Mw�┈;.��+r��0��1����$g�hn��ilf�ʵ����E�Ղ�9)ΜB�$�;�������P5s5-�Y�r��>6l_��h������|����ݭ�������kH�\�fEOO]���	XR���?�vZhl��m����A�v
��Y�._?�s�����4����O/��ߣ�*Y��.�總���G��&�)�rv-o�@AR�!����Jڠf�Y{���"��^���ɧ�^&G�
�'n��E
�g| `��/�z��[C�iU��	�h4_f*���~��
�IKKwttX���ި�a�ͣ���&1&���Ma��V~��J���Y?��p�;��_��!�Ɏ��?e�Ҟی�V��
*O\�-�·�g���Pj8���U$��l�I��������jyz��
\-��������5 C:O���D��?e�*�NQ�)��T+(�G���:�SÕ
 I���!^�&s�H�\�g�ΗN?�T^vƸ)Y������o���p��E,��5��$�B�ӟ�f����<Q���̩iq~i������f�O
[x��bF��׆LE�w^�_g�ޝ]��Ib�X�v�����w�S�͍�AI9		5�����u�r~�'�RR�cIl���J���3�V'᠇\>���k�M�N(��d�,��ղ	��N��Zط��b�=�$�/��q︽>�fƾ���qIh����j�G��+�:ϔ3%SS�����ui�F��&f��I�G�-�U�!����v��j3�CMx�����O	�*����;}��?V��5�&�$y{d�C�,c���h@|t��ށcԢ��K>Wl�'т��|��˓�����"�c�c��S�_N�4o��1�xgdFD�s����D�ek|1�.�s�$�����x16�
�YB��&����^�LFi�[��y��������Zc�}^(��Ϸ�CK|F�?���}v˯����Q����ɔ��?̦Kk�&�ʿ�rۚ>e Վ�Xb�"Q���n&�>288O� ��gV���<l��=�Q�������/󟁏�Z�+9m!��h���X�0W"}M���e��b�=�wx}�3���8�B��4�8���F�e����S	��hD�^«tq��Yd�7�R�/�J,-,�X�(&}W�V�*k�q�����p7����}%=US�t.�3��Ej��c�a��	���E��q�0���
�}����Z��K#�x\��.�-�F�l�I��m{����2�Cäwۉ��l����3�9 �����O��~�E����_"��S�j���m^�Z�iU����;>\W�O�l�0a?a;�ȸ����Ѣ�w4���7ӈ��>d��շ+T�f�K>XKqnn�吣�?C縭/r��/��~�/�u�mD��`�x��&ls-g����p�]�]�W;Ad�;w�&��VN!�p�v�u0v�n�6�v�^x0s�)�vi������ZV�+�_}$'Ff�up|�+U��ĤU5��V3*�䣋�
�#��M~^��Jj��A�^A��Ք��x?2ئ���R��������`���92#]�KH��z�B���W�'�Eh�C����)
f�.:��0�0�{@h�Cv_*���G���6B�<5+�h�'�:�ڥs����.��wΧsP(�J0e�=;���g�n�1�N�K��W+�,X�������ڸ�D�&���s�R�;!38��[u����Ʀ�}
��O0\����O���F��N�N������sw'H�A�d��_4�g�A�x�0��.Vk�ᆱ�Q���l��4{��9��y�NzT!cj�8��A���cB=�<B��I�Hz�
9�� o�ѕ��|ҕ#�&r,���n�4ٚg � t}�p�|$�c��BF�ĊXJf$9"O�9�y?&��?���H9�TZ۟�U��7�9yD�o��f�<qЅ:���@��ha���������0���mٟ��M�Ȗ���"\��f�)� ��>��y:U 6��	�5)�vB�[R便����E�i����D��+���쑊wo�3����.b��gӝ�>������4 z�Vh��\pTS��mKJ$�kV>��qc�R�u���S!�G�����(%�l�z�>[�G�y���-[�~�]jv�K������(0K~R���)�K�E�K�I��ů�J�ٔ�d����E&m���a�!o�f�����}aڥo4�֜kM�2Q]�\,��g��%��`v���b��g�i��K�۵ɤ+-�[��@W���P�˙o��!Yv���e�D�^��UN}�+/.�#��V&z┏�hSf���%��(��~Q��Q�z=ᗧ�>�������{�TO�Ҡ�S�+)቙?\�RyZ����h��&q�F���΃!�	�Xt��%::ENU������l3�0�\3;�R؀ ��?cSS>}�ks�����l��L��"�F�pJ�����u�U[V֑�wx>��C�!���G��A�g1uO$�V�����BIM(l�8�YTd�ՙ{�f�=Hk�fqN�����4��O�_���eNH�+ܔ��蛾�[����c�R'+������P��h�d�C��c�7XWJvҭSQ�N���jO�yn�{#� �1�]��vL���q�8��ơP����b��iemaዋ�q�#�^-��wEy�A���	噣��}�����5����$۶��@__��\��&o%�-�8>�]�����@�x7�$dl�Ί�%N����2�A����4b��9�	���B��^*��o7r�V�
��6�52՝�?�[�Тġ��9�G)�k,�s��#�[�tF��܅g=?�$9��ފ/,o1{F�+���p0WzZ�T��$=�Io(��9��:�FKk����0�{?��<�X�ƽ&JUg`�`���9	��{ł�%�阗]���=:�W�E�UP�y�o�2����Z
�(��J��ީ~%�z���y�0�k�qk�^��%eee�߼�9w����޻¥Q����5�*<�1�!��*�
�,/�| ��%��bOఁ�(��OQ����O���������#��E��g�̽�&z{:�41o��k��t���i]3���8��军�h|��#�z��%�J Hx  `t�43�oб=�A��6��-���.�&���~dĴXl#򰿶�ۣ�"�Ue ����:	e�}�ކ*-u(�bGD 𧅔�^��Ƅd����6!�s�O����ӌ�5��w�aN�on��YYY���-�����`?|ػ[�5��k�b�5���(T6��+G�0K
��g�n�/��>1�Zx%�2@�����OQT5?Dx(+���<b�TTO��E�6���\�a��"I��R��O�*���v�>�R(���VSQ|	����p�G۝�j�6l���,V�*�\H�Q2l����#~T���~���H��Ė�J�������c22 '�𳦦2F4ԱXli)H���9`��H_J.�p=�����`��ߺs��J\:�A<��(a��a��p��H��謶(�h�����*��q;�:F{4.w�+dٿޝ�d�+JR�Ւ�Ʀ���b�}9u��Wۯj��u]�R�B��/m"<Ϯ��k����wrF��]D\�IJp�5�{G��Jpn7iq�m	���Ղ����]�Ο�|$��5��;O�]uԇ�M���"�]�"ð��MI)���õ.Y����ۛrJ� q�B!ȒRtG�� �^��DQ��q߇%�~���Z�l{���-���/1
��W�I}�R˙.�{�·	��-i�<�}��J?�� O\� ���,��{8ώ�ߓ1ns�8��X��-�<m���u���M���l�¤#��G�M7L�������d�ӯ��>dt���2������_��/�#"gI��KR��
��r=�3����1��R���h��`�t:���87w'�%����������ru���%r�c}�!\`	P��q���	.w���������utt�e����d�����7�ha�C���c�f��0}��hz/>u�п|�g�|�GX�m��AX-Do��y|n���1�_���=f5Ǵ��!�J�NF0-��%b�/�bb�q�[R%�����1_�u���Ŏ��V����Թ�����v_�B����Z���x��8j�5'Gǻ��I��u���r���^m������b�<�T_��h�kO�)|Qy�U��=b���F��_��1�M�<�|,�֪���"^9�����
�n8�G�$hX#�������,�������WI�����LE�ᆦ#b�h�I"�����Ŵ��A�p-��z�Z�s�����ڇI�PC�~B�!�(~#�S��}U�2S��<��0�Y���%�ay@�AL%g�U�I�=�Go��W�%�7�R���o�p��RX�����3��R�l+�>�w����H�;�����K/n���i�<����Ǐ�ls~�������U�d��g��κ�oW4�-f��c��ڼX��\��6����1�����~=�{^ߠ�B�~\� D�6֌�B.֌m�P��\e�O�EE��~�������;��::�C9dπ�&�Y����߭���v<Uc�B�f�=��.e�&|���D�Wӷ��D(���kE�Q��i[�������q�k$6��<��Ic<%ǕHe}��כ��ݳ������{�1�W)���4���<Y"�=��:�Ҵ���n�@a��[5x���P��*�	����'�±�pzIa}�:a$u��RE6��dUo�r�M���A��'B�G6M�W�%��/F���{�t0�͚��@;b�������LTaV��Ly�Ρ��Hedf�K�V��Ί4��C��##�롻C\��W ��H`p�����57#h�E���:�Ni�UoT�����a0�*�^j��k�]׈��G��2��
�X����=����e9(��d��!Z~�?���_�E�5>���.##��/W"��]�M�/�*��U#�Țo�Tҋ*�*���[$/�E��$}8rA4C�G�[h���
������r���uM�/3��V�R�\1�[��/��3��}:���e�o��ga�׻(3��x��}WU��O�+�LnUL�cRXY���C�G�]���M&�0��Wbv�Q���Ӆ}�٭Ě�Jg���o���~B����ۖ��m /��6�F#?���~����C� ���"� �c\�/��=�]
�~Fx}8"P,+�rV|.3��@�)�y=����|�^QI�;��h�J�S�����l�A;$��!��B_S�+쾚��{匴@�M�!���t��v��n|���!<ի���J�a�Dʾ$����/��YV�����K3�ctf.���Ml(�C��93Be��C͊A=a=}J�Mau����R�b̷�/��E��ӵ�T�OW���79�����Ɣ�/����t��x�r�'[?��z|��e�������.ן��f�ӗ1��Ӈ}G�),r_�<-��󍵜���;���F��l�?!/MjvO'����ş�f�	�#�1�k�-�)����P"����V~�����(0�@f�7���*k��!~�8J�9U�#Z�w���P}���68Q�������}D|0�]����k�����۾�K�O��k��y50���]q@y����i�m���~4 �Â�X�����g���I����K�%�)YB���V��1��zR��$$(�=Z�n��m��}���SG�#;'��c3��o0H��5��:i錢��?%��Q���g�����5�{v��tI(E,�:|�$2A![�gQF���d�1���}���|�u>�{o��>@h�7��.j�g��x�m�rDW��<�<J�5l\������.���g��pS*E}J/BmvW��İ		s�>�]��]^ؽ���!x�n	�|����N�����hX�<��zӼ��
� W�ձoՔs��X�U�}/��/�M��/ϴ!FK�@�8�5��A�F��d�R�@A2"��Gu�}td�4�/���Gۨ\ݞ.캤����Ք���ϵ���s����I,��c����鿝�Å]TÒ�4��h�c\9D;��E/��!#�Z�DF�=q��*  �B)�}(�9��;����.�����^���T�1qZ���F�����*:���vi���`JV��3�A�0�G�8cutWT�r���!���j�8�6��H
;�2��p�7!��Z77�mX�E�F��Z�ќ~��|�\�U�Ȩx����^���҉�A@WZ|]�D�Z�@��k݈q;sd�])��Ӭ$�����l�U�-2�	*��6})8{�T��ʕ��3�x/�&���uR�Б[��V��u�o�,��c�#`��d�|�#~��u�ڷ�zwp���W���[_$�����;��;���j%�� �ݢn֝�/Ě�ԧ�S��pq��:l��*�^H<�b����������z�vf����qǢZT���=	�)��*<��T�����<��^���g2�<���Fy/ڗe�� +��/�(�N}0�ٳ�X�4�LKէʲ�g��.�X� ��Q��n����1�N����[_��g�ķ��H{bzf^:8㣺�O��}S}������TYX��I�2&���!|qk��T�}�F�̺��Ȑ������y�)�B�������"���k�����K����n�`�����Yl��`������vw{���O�Ə���J�,4?���Ȧ�_z#;^�'��U�Q+u��+��ͧ�Uz>�˩�����m5~����j㴵�/C4�E��#vk��	�~�[� ˄��*3A�P(���֪�uyġk7�Eq�L,̆PQ�d�����yR�g�c%��i('�2���JfI�6~A3��L�s�t���C.�����Vc��á�å�A\�KHTo�7���JaZ�v0��
��j�tD��� �kT�u��:%ܷ&V��GU���J��-:%RkKr]Rn�O-nrɜ����]Շ����^P�ō����|9��4#�*%�3X�K��qZ|
x���fS�I�|� <fi�g�UX�N:�J���J��^�1��t�,	�p�%`���Qz����C�ţ0k?tl�����5HN�m���N3L(0�b)�||��Lf�,�R:��D�m�-���*ҕ�R�j�D��(��zI��O�Ȯ��w�9��I���a8�E����WcG�6��Ñ�e*鉖z�ϐ���M49�EՐ�������5T���r9x�������^��K/���]��3o�X
h�8H����X�ìLL�ݸ�Ҹ2�-�q��&�T�9�`0/l���8�G.�d��t�����C�����������9gmHb�����k�u��y�5!o;�\��e�{�_���yJ$��P��U���T�"�GW终�H��~����˭�>�y8��R!O�3%���~̬�oI�l�Q����B?p�����t9[4�v��N���
��ɡw%Ы��%� q��'E>����n�E��bwg�)�O$��l���7
�]�o ���������V��"(�g��g���_��O��/U�՗��*Qz}�&������o3��Tޢ�¢�<SÏ�a�B+f,�D�e�� ��	��_~���6?��7�g2�j�N�ў��x���?��N�n�dV*V�?�����h�R���P�R�|ߋ*���P��4,.�`�z񑗲�>��	�
����i����V�TH�#ձ���pG���$�})���XF�(*�N��[C�m��G\K�$�w0챈���Hl4�Y��:�vk�����������y���=<�f��9;J��fdd���K�sr�Z����'Jh�ػ�=��߭���j_2DXv�Պht�_�䁱�K-*�J�/��1�Qhv�P#�`L�>i��Е���a�U
P�k�GX9��a�\�*N�&S3���A�����&�M�QMgKW$*�j<Pj2<}�y�r��e�����d?�h�(CW���B|��芜�𛍃���w��BK��!��®�3�����'��w��"������t�>⧮�RG{���W�����|�G|�I���[��y����:����S����|l���H�}K��b�oy�O�uղ4Xqaqa�x����uR��j���k �ci1��o��m��;H��;8zg�..�V�ŨJ�3C*26<��DԼ�����͹�|��jN�%(*����0���7}�ޝHe��|
3�=R{vX+�Z����2!D:����c¯�<�b�⒌?k��I.gA��I��NS �؟����H�fr��0@��R�I���ɢ��� �g�Ў��m��vv	@�>�"N y|���	����YNL_
�"����Μ-]ne� �%rg��;:C�/�.�E�Y��j+�0�t.��?˒⒢��O?vV�m��戋_E������0ueT;t���y�Z~��6E�L�ZΧ��b$7je�x��z����4k,��H��e�)����S\�=2�y�d'�ΣP���	گ��щRvp|�Nd"������J���"-��Y�v���9#}nb��^M�El��b�"���"�!!-qV���X�><<��񍈈ptt���

�cLV�هfj�XI�"I�:N^|2��o�SW�'����أ���5Q�S��H�j^ѻo�uJ-�V��7&y�uԩ��R�O橠ʨ��4�˙�zP #�D*�M3H3��x���'��{8p% �&���H$�t�h�ndI%���������`w<7 �`tl���UPBz�v��p�/~�!!�K���Js��A�s~�*CQ#m����۳<RE(ދ��<�zd�3��.�32�m�`oґ5P� �,��5,**�B9�������aeH��iǋ���D�de-�iKB/7��A�M�˥�~��r��ڬ�x�ZNd�<z���8,��)v��3�3��J��rD�-��C���w�ѣ���x�&6F��z�O ���sU�����k��
[Bf�?�}�mD��`�1�;�g���Wc���5��FϨ��=�]>�Ў����Me4�D�q�%No=>���*ڤ*��c����3$��&�Qk��D���c�d�+��C�|2q4��,w�X,�Yț��L�݇~�{N\��q#�p�� z�]o��T�c�	V�h0H��}��H���;gd��[<�ԩ��K�Y�6���������1�J˄n>�YV֒���L����%���'K尌�(h���)�)��J��⎖��֓���[�!/�!}�5�J
�:�����v�Fjҏ{���l2R�"�{�&,�O\��r��C���:R������t{����:����Cf*���,�Zr��$i�Q
C`
 e�p0��5���@��Bܮ�;���
�#³YhcW\��C�cee%P��7N���*k�C��6Q{��6I��}�%���7�^+�Ƶk��uF���a��7��?<�n&X�n9ɴ��� �Vk������z��|�l�x�ɦ�x_
�c�|-����*z�n�,*x;1u(L���jh�I����Џ�[�D%"{��2��"Ǭ��*����|�qOۅ[�V��j���߂ja�O��y�����S��'��~~HG�Hb�k=��d���]�G�?�62�����B�������ت�S鱇A�MF�oϣi;Bԥ�0!/����v�}6K��h4���/pQ+���eW��:����ϭZK��t.h*!��[�Pԟ
�L�/]��m�R����)wK������>c����-kHW�cOhY58B�A��3)�%���s�+y5�����F!�gD����)ɑ0̅�v�@4�)�jW^B�|GQiN�`^���X�"��>����;x�2\U������}yt��ɼ`��#'�j �:�B
�S�Lo�d�2��削�>�**QR,:�vlӷ�j���#�V���%���D)�=���@���O��%�L�9�]�Kn�L<6�r|������ى��gA(,Mk�h�ś�xڭ������yO�:`H��t�=x���a+X��x�d��z�Z��� � X9���9��H)�
�Z���H@��OQ}��@�/�m	�^���Wl#��,��'�]Ĵ�Z���ǘ��J���<B�w߅�!/.����Z����ꪍ\�o���۩���U�p�|�N˅�N TUU�0I���I϶��\9 �j��ۯ��*�7_7��!������V��k�2ۋ�H-�g����G,ԣ?-.���L��p�K�kj6g5l5�O�.*�}�N�P�Q�R������������`��*��i������2`�Y����v��9���f��|�
��E�K��*��Z�u?���fɇ�N�wu����S�g��lC< �4��N��_b��S���@�]u�'�S�H������'��L�e��0�ø�8,hS*�R�H�T���L���p����^�FKͮ��T�ǳ����cb����l�4찘n���!-~�✿�}[q�z��al���|��5��-f��Þ��,E.��>���H�O�q�ט'��xI@q,03|"�����1����̋�|���c��-�1^��]qr�ϻ��#�� �#�m? G��C�:���*����c��à��I[A�~!�YSb��.���t�f!�~~��C��Qe���B�O�w;��|[ѯ5�y|}��P@.���K̡=�}����ubQ4ԗCxi�Uˑ�����v��,��E��.E�������\\\5ER�bZ~�u�J������3���'3��>0����X?��DkM�)���ݎ_�nl�q+��-I:�G��L&�`�%�n�0s���#f'Ȓ� ��eE�Ĵ������gA3	�F�G!��\�^�mH~�$.�}�n��S��G�֬g�-W��JJb�Q��γ��:�,��Lð�R��j u��y#}!V�/��t���7����W�q���
��2���LF����o�
�� ��e� ��IV��9�e��pR8���m2tr���o�<LX�tRMڨo��b�H�_#<�)�8��$.}�))%��	k�v��R���"�q��^���:S�Y稍�ׇ�( G)Zn[����Y��W�����_	U��W�[�=࠺�`��Vy��iJ1t=�8[��!^���D0�FT�GF�:�rPM��OӳG4����q��Ab��v���	��O�O�t����g����I9��O#�u����Y�@���>;&�l�x��i�H�my֘F��B�׹�o� ��PbۿI�f�����^*��~�J���pڗ�q(Ò���~`�9��p���1y:�L�?T'�Mb�f�6�};4��t�A*�0��!bY��:4a5"m�
N��\�� ��>��b�Xk�|·��/ʣ��{>U3^�:��ֿ�����v�<��hKEF0D��Pt�� ��c�K�j}�{ĀtJ3���)�[ڤz-��>K��1A1����q��N���p��۽�C۴�����Z��,��zVP�=H?H,��e��(���������҅�9OJ��"�^�- ߭��wтЫJ?���t?��o��M���W�G�<��O�d�}�
d��5��G��>��=�j/��W�J,�B9l�1.�Oa}��~J���b�Dp)������@!�WB,�K��R�B��Y�̈b( ��%j`VK������CsrV9���螉j�OϜ�����U71ii�����2I�����`?��Z��d�(�@��3�'=Wa�C?8�w��=���[
�JI�@���2�v/5�{�I�=a䤒�{��2e��/�nH�h�'/�ܨ����RԮFn�Lǉ�^5��sj�0����$��K2\e����͓w�T=Ww�Y�i�����M%����X��?J�K��>�ě{*]bI�+��%E�W����!�l�H��W�P�6-2��4�2@E��y��vZ5�rJW���*�^	LUJb15~��R>�U~��u/a��̶��ʑ"9�z{�U� ��@�bU�Ti��l&X�#�����<�NS��c���q`��w���� uny�$�����dwp0��~~o;u
HMC� �?��U=�h�U��f�O���ϛ�ĆA/��׏Tl�FsA�TZ���o��]�<�NS4k��]�e��!�I>��'Vx���|P^8�`��-h�\�o��E̗<� |'���rk���j�+$l�Dy"Of...p9���i��Oa�$�!�
�d�|�\��~��2!hqKLu&�͕(�;� |歝��dH����ɩ�@�����T�ͣԲ��$vjh���5�:�144H�E@���J��͆�c�<�t il<iQK��Π�Q��[_�Y�q%a�f.�FDsbμ�M&��V�,L�k k]�Ȧz�`c-�c��O��k7Mi�Z�S��XY�t^<��^��2R�>��)��%sٗFc*l�{���E�I�HH�_��&�;��f��nҶ��>�X�{�+	�l�RO�NDN>��QllĭzO��4U$�D/�0��5�/!��-'R�~�d�S�Y�v~��}��f��R~{�6^Y���dj��%fĵD��� >D'uwfL����X`��셢�&��qjcv_v_����U���vuu��>�]�?�E���D��L��.���K7��'c��rl�f]A��0��³��(/���賟���x�o1�o����?�Y7K_O}٬�Zg��3�O�{������O�+M=C����;�ۼ�!|�!L@Z&>�����v�#�{��ʹ��KU��Y�8�&3�������2e���\���e��S=˧4�e�$<g���b �ɥ���b3 @��X�9N$J�=��G	�hu�aq5'�5�@*3?N�xy�_ ,B �}Y��P��l����&��ϖC/��ߴv8��~%A�|�H�5��Ʒ����b�S�����t�\���=��T�t�mX�	�Ն�B`L'�s�WmE�"��9�s�U�q��ؙ�e1n�e;0��/�Nؽ5@@�~]�� SO�}�ٚ�(d��s&|� x ੠���|l�ϳ?u�ʿ`b�!Y�Î��੢��o6ޫ�J��"P9�׉��j��Q��sdG��<�
��<��`\+���^�'u��h�N_nll|�[_�6�8��x��[�we�?$�����+m���%ʩ���ЉDO��%]{��a�I��l+G� O��	���2�����������[�+�幃$KS��_{��E�$��+eQI�Bu��H�o��R��"�,2E��w���N^�>2�Ex/5�nO�d�Du~�,��%��z�����GGU�����c`R�J�Sgj�_�w���_��y��3�a ��~��ٴ��C���A���J4Z�+�U�UU� J������r�^�$6�0+O(C��zP��7��3����6/KMS����C�}�Y����Y�֘sǅ��3	B=���q�O��ʣ�ĒB�=ڂ�����~��ϼ�'���l�P�%��Q��å�:	���oɻx�8d}���Q|��G�W)s�6�OL�$H�bm=Z�4��o|N����na�Et� �@U�pe$��$I��\���fT��v��lhJb�Wˀ  �ʁ������t<�	!TU5�N�>=�!:��ѨA��ϟ/�]��R�L��	efVk9mB���F��%UP2C�
YoX3G�@D��@ڂ4�2�&���F�֭�v* ���MZBUD;TUT��R��4Y4:g��d�RJ�����8�j�ٹ�h4�����LkVav�^���Z��W��Y<m�3;�e�~qk?�F6[y�6[-�$"�QJU.}��ӣ ��y	������B��i��@!�hį��lR�d� ��Zlɏat͢�W�0��Q"xc[��V�=0j����2o9�m��Ì��ݴ��H|��'SL�
F�ÒP��{�5U�[t���.|�u��3��J"Z�݈�!����މ��%��L�A��"1�h�����B�]�� ���>��|���Y)5��=��)��V}L �$�ߓ��K>���%:��_��^�Eӹ��[�_{�R��]��L������;���������U������]��ɋo<
��Ѓ�(�k*7�=�HUC�b옐���k�d�=����r>�N�H��u�P�oj�-DH)E$b�|][�[Q�놘B붭E���:5�u�ŧV�ժ]Q�4f�U�9gd��jU��Un�^�V���pggGD���δ~�CB�\��[��_�-u�T��&��Hr���."��M���޴}��ovq�����4���Z7v3�@�Ɉ��wm0�8�$*UU�F#�S��d=/�+Qm��.���!13����$"�lo�x� ���P�ju�E�~���{��:��ʛ���=ԼD��H�m��e7������"�H��ew@ FbI���I�֮DT�<2�%c� ~fǜ0i�Wjadj�O� �9C�9����$0���j�XΛ��h�4u�A@��	�)%"L�$EQ����G5�o�$��f�������_�#����9_U~v~����x��/������mۓ'USIJ��' �$�,)���6�UAf� %q�`.P�,Ki��H%�T�dZؼ! 0�j	U!f�>x(��ٴ�	�%�!� �9�b��1�VUe�fH
��C�ʩ�FM��� D5��Iz��t	V����2b���BD�h,|"L�6S�̘l����#��ĀZ�-&��¨�VQ�m�D����]Y�Z,`��@ЬCY�N3�3���y⩪Hqݮcy��e���D���Vo�q��_3����i���\� �׆(o��k����P�o����)w���k|n����%��"����O�c��ߋ
�H�܂y�q�Iu�C��+-�D��	� �e���*I��$	9�D�5�B.��z-�`~�*'�@3�cH"�4kĵ9��Z$�S�lDZ<,f�QT��e���n�6DDf��0��0�| i��� ie��oh{�?!"�������?������믽�Z���w���������?�/�$��0���m�_�i� ��ٛ2�'�W�f#���vm��1k����V]�bbk���������A�"L-��MQ�j���i0�S� #J꺖 ��ж��TU�/撤��w�mW�z4���Y-��r���3�cL��� 8ݙVޯ����|�^1��r���L�[���Djy�4Xk�m�l'�r�M^��W���q����u�w�S�
̮�jk�H1FC�L����*"f����cV��D�k���nh�γ�� �$J=�H�l�5VӍ� bJ�{a�d�����S�W+"r�Kp�pZ�l� )�:$�~3`]�U<u�D %����o;��t��t��D*����c���+�����j=#�M��x)�����X��6��x� ���ZN�{�L1��r�Z.�뵚L���mk$c�bD& GĤ�9�k���3x�^���$�!�zq~~q~� � �5v�\��bj�>H"�o���s�� l|$�ɔ{u0=�z�X٥/k�X�f�T�p3�:(:�H�M�BD� i#q�n�u�T�8��P��AV]Pfr���\ň�S��`�/�1E��0Ѩn���]�)�
]�V�uu]���8��q��!��W��;E�N�Y��]hq��eyڎ(�L�	�Uc�]%� )!�!y��Dp�t6�ΡtqA5��Xa���H��I*�WU7IBp�5M�}�H�\�u]�=�š�y�"�hY����!��b��-�xZS`�!����e@���t�s�ٔ�im�p��@_wdi�i���a���e�;��z0���a@!@O��M㢌�"��B &b�=9J!��:�[����!iF#U5o�m�6�G٠o�,�c�yh��-j��&F��וq�o??ĥ�!v]�X,��ݿ���������ʏ�Z�sՕ�����M#�������
�ie���R�\XVE$��� 0�u6�dˤ��{�(*_�cD5�H�c��c�v���K]�1���Qӌ �yUK����c0#9�ϙ�G?��ѝ;��ӧO�x�W_{��O>����_~�қo�yvv��GTU��o �{���o��z�4}��j��w���G�>������x|��W^y��駟~������Wu6�}��Gm�6rPqh��_3=���i?�&�[O� 3�P�����f˦�HekJ�6U��0p�DR��2	%�(*�D�P�@A$�p�!���8v&�j�.l,���j�IUʃk/� d�QǙ� �l��@�<"�QF��J��le�ɒ��u���y����Go�_*�ߩ ��Ut��M�x��`�P�5M��D�0�Kf�!�!)�˰�sKM��Ye8��#l�{m���b��U���'b��$�0���q]��X�u�����3������ԅ����}���5-o��e| ��*�c�I�)EP�u� �Č� Y4,{� 
�!���f#���5�4C� ��w��$A��!;!ژ��r�P�]��t����ی�R���N'�V�r�tB�$���QE�:溮�f�v]�,���}J1��u]3jvFf6f�&�1���H}�K�����|*n%X3���ߨl�(m$��i��l���{��g��fM�B
�諪��WUe��@T�jΛ+�T��5r@ɑn!t�����*�#U54���M�^zm���%$�P&�/���Ǖ&��Yu���2!�ڀ�eW��o���c迼#����th��j�)E�{BH)10d�CV5 }: `i� 8�뺞������yA������t�-0Wː��׆R&\��i�]P��q�I}�o?^�Ԝ<Q�u���?��������������v�U �*)UU����o���O��?�/����o�j�02WSje��s����5)�wΥ�s߈�ДDU���Δ��C_�*Y�A�m�x��$I��v������A�Y�׈xxp��_-�$�Ν;)��|1���/?Z��w߃�j5��9<8��Ï�����×=��/��t���o�����0�^�����O?���Z��釬߆�����Ch�y��y/��F�/��f��?P("�7ڭ��60�7L�.K@޻����eb�'"�)d&Rͺ �HD���9�(t��Q�F $�z��=asu��QM�L�o�2��l�p(͏T�tm�fGLˣG!�2>�/�M��f��?+gY�d���M�W P@Ѥ��Q�t�W
��D�>��6ps�-#�T�����]��V��+���q���"#0P)��ߩ ����z�'�q�4u]3sa�^����=a����;؈�138���w]��@[b&n����5)����3�J+�X*)r>�S�v�u8�[o Q����%I��#� ������<8v�X�V���
U�ZHI6��}!?bJ��:D��{�bH)&g����L�z�ځ *OU�1%� �)��뺮�9�d p��㔒cf&v� K�w�-A@���@n_�ڻz���3m���xb��7�10U@S{�񊖬��x����b���L�����A�9���9��$���%���3KFt�f��(�Sh�uѤ�J�FKO�~����ZbR"��&����'�	�x��1�5)ڨ��~m\{���
���YÌ����z��g�E�5lj�Y.�?���hvJKB��|�_/���3iJ�y�y}�č���k+b�}�;�2�b�#.I~��\fY������_T�O��3�e�s1��r����;��;��w�ɛo�ѵ��U&t�$�.�n�S������.�»�bH���\���(��VUB&b�S�CY��+�SJ!$�*�R�"D $f�\J�t7��jgU�ڪ���^�0��F!�6�~�٧���;I�ɓ'��z�X0�/~�ӟ^\\쌧����o�ݶ-���{�}��.t��������ONN��N��:;=}���N^�ؙ�c�|����e�Xh���63pk6�^ YJ2w�͠D¬;��ޫ4
����=�P�e�{z�v6�AzoESL�x���$�lGs윧+��6����1[z'+<�Hiq����pR��%�e8�>^���<�3���H�X�kj�/���L�D���ݜ��r.�a" JIb� Ztn�r^��-��n2f�wx  ���14�h��e3����	R�NX�@򖉀 ����D ��kd����0x� m�^\\�`ݦRq�[�»��*�%�bHA����9@ @�e�UU�J�%%#O�]�*��Bv��:&Xݷ"��̥���B�¯-��H��o�E�7ߴ�#�H� B��;f�焪�T�dˬ�DU
���-i.!�R���H��.����;������F�D�̀�u�
3�������m״	�'��R�"z��vlt�¬�����\�7�ZY�6۠��ιd@ĕ�<��! ��l��DB�=i�d9�� ��7>2�f�xM1�]B�U]5���}�M��d���ֲ���_e0L��D_�]��D�ъ�m��h���Ө�kR�$���̦A�:�uO�� �ub(�����<�i��n%�o\c�[�X���������&�+#!!9�*�{�P�1���&�5��d溮�� �\����n{9�n�{(0��Wp�E�Ř9>�=RF�W\�+'�s ��g��i
Ɉ��b2��{�����������_[/�j�T�9|���py����ݿ�� ��������{�.����8}�d(�+�`S(3Ɯ��UPU��ƛ��Ő��L�e�I5��X,&w&u]l���pY�0t�&����t�d�HHT1�u������fO����"ryy���xxxvv>���f���cl����ݿ7jF����`�ѣ��h4��&���*DBt��f4jۖ٩�U�\�-C?�:;��s��`�m$�`�������Cl���;Aqo0�"K�X���2���/6�-RU2@�p*bq���H�����d1�mk�.�A�U�m[���$,��?��YU,q�P ����|�]�d�;l�a�Jd�:�/�,�f�[���������L���� W.ߛ)}� r�)!(i���d,�)Y a���vww��S"캮�k�8G�:I��˄]��!`����:�IM� ]O) B �j��%��"�#�͛� H]U�=I�׀)7o%�لS�
������VA���H @M�G�v��3�T2�n�;E������㦜��͌-�=2QQk6\39�ͭ�\Ldk�l	T������ �Hr\pMDDB�"O���\U�L�b���0�e`u�/DB귫l�7U��v���\&��"��B�XH��O��mD�2~�u�DD��V�n�w�k,phj���@!�B`�ι�Ā[��������Jy��F�q� ��#����`���&�E�m��M�^�~�Xz�w��W����p�t�g�<�ṗ������6K��d�п�m"�xa���"�y�e>`� ]�um׮��CK�h%�u]�u1%@!ꦩ�_����М�(�?@�I%?���4�A�a�Etˣ�B���zow�����������}�R�b}k�
��$)
�b!�{�����;\�?����������z��jѢ�~��Q8 �����#""����8U5�x�4�Y �l�aLڮ[f��ۻ������2�:����]!F1�'D�L&��k��K/��X,NOO_y�����'?��ϟ={��������裏�??�{��_����ɋO>�dwo�o��o��/����o���?xp9���]�����W_���>���^��_�����~�Q��n���- < ��|�KZ@�oIv�k�m�A�R�Y�I�zdS����3��=K|1�|�%�j�d:k>c
!jF4�X/�.t)Fʹ.)�>׍��w4�V @�����w��޳��:S�c��4���۱��o��c\t`�˫�{JzU5�U�r�+ςWND�c���a��	B{uĀ ��C喣G�T��W�\U�9����+��P�� QD���^��E�` [�u)ED�Lf.�M<9v��&��3M�4����_���L����>s�
�j��D$�0<��E�:�j|[ؤ�O�m��q.*��Dд����W� �L՚ʨ�^��xɛ-�̀}>�Ric�&INQ �
RC�uc�Ns���aNY�s�
yas"r��"�lw�}��楖����nfr��@!�����<Ӏ�˫.�
D4�/q.+ �m�����]T���=����Pb�,��))f��t+����N�i��s]��y  ���C/mp������p��@��S�6� 8JT$�U�
���c�_\i�s۞t�������{��m���`��	mYjV����V`"GD��j������ ��SL	��{Զ���x�]/%	"#��XOK�\����6
z�[���-hF����j�>�<�o���a9J�����.Ii2�����������_K�R@r�ɚ5�d��d��eO��w�vո������cI��l�T`�����f( QTS�z#����r��E� *��ܷ2SUǒR���Q�Rj۶�����d<�͞>{�Z�.f���d����_{���?x�����g�����������ԅ;����[�5��?��?~���o���y��ܽ{�~��f��?�۽ݽ���ߞN����?�'?��O^y�������k������O�>U��]�uS�� , &8H`Z��f�D�R!���7�(�>���P �-�
�� ���d�6�齇� S*5�"9��bLTe�QU�z3�P�*0|�c��W~(��)��ݚ5 x�KU� }p�;9|'��e����_�@@�rd�+�r�9�f��7�)��[D��`2_K�CepF�l2p��T��`� ��!2�1$+y�ؖ��,�
��3��2;GQ�]HD[������p2[6����RUcX:�T5����d�KII4��]�����k[`?�W�׌&����}�H�iOm�5)y�\?ڿ���s�QRI�F.�%Bk�n�E&M��a�C�.x�%���fJ�K��-��yq1Z�:�H���Jb��SQ�L�Y`�A�?�*$I�ȊX��0�aE��qk�@I��SUP�՚}p>�}h6#�H�]�v/<pe��e��&�9������.u���Ȭ��FS	o��[*�s�����b]A�+��&9��v�Z��[Y<ƒ,��r=�.-&��Kn=,C����u�S�(���tCu��huH6�b@��t��o=�_�%��%��b2�1��-;�VR`ʞ�.�]�y�E�C��m�a�u!t]��P�h�;#��ܳf��7�ٸ1�"J�Ph��o���\-b������9�^�~����?����~���r5jFw�=ד��Q��������'�O��'��Ν;�������|�X�7`��֎KS^��$�zϒ��F�4�T��:vD�\,S��r�/���2;QQA����CL����Ν#f�1��Q!�T�V�1(�z���f�Ւ� e�Z�d:m&c �����x�R"ǯ������>��p��x�4�x<�{��믿���"�?z�{��k@؝N��߿?7�"�ij3���Ñ�gPs�&���c�t�ڄ�NWb�\�f�K5d��	�����������ED���,�O]��;/I����D	�|Bt�!�m�=@p���o�(�1�¥��~�@Y����^��@
z�ȗ��*Vڍ�-�:��;B��m��nC�T�%�����,֗�r�Q�:�8�*�5.�w��TU�XD�1K��%&3�D)ƶmW�e����r�X4M�W�齷Z@@��b���oێ���8&�()��,�~���64�P���E���I��
W�����Ѿ��t0�g %T�Ac$4H$k���gb�fm���J|-�c�|�������,=���B�"�x<��@s�h H�L$��6.�x<&$���Q� �T�@	)�DP��*B!H_lX�cP�d��v�*���x�-G��Qю״iw�����M(�`�;�w���`�B���̓�(��y �Sɼ�3i)ݰ��U�3�����U嘷��n��m���"�Ͻ���p-�}����3n�vˁ U1��T&)��t2�J9��ZD�  ����sۆd�������{m�����Oo=;�����(�����_���J������M��;�h7��	Ab�ԍ����uU,�T4���;faB��h�3���s�ј��U~0��+ꍷ4to�*7����a��$D�]Ym��\ǭѝ�GYc�#�����$H�y�#��.�;;;���������?�O�pzv����w������]]) %�&�ӌ�����������v&��4#����P3ߞ���	�E�d�&"Ws�n!q�v�ڶ]�ր��@D�*b���%�<E���j�꺰���^��U�
������|�4SL��1��k��?������/�Ǔw�y'�������/��W�����O�l�j��������/���ӓ��o��������'��/~?�8��<;;���_��?Z�]���������ދ1�vs�M��U�7Ύow��~[1-PS�o�Ʒ�'XX�jDIN(b}��q��M� 9b�v�Bık%F�4�7D ����?xo_�0��|O7���/�VD���)*����=o,[�[� �l�0[��7�Yr��j'�\�eJ���}T�6����G�6�py��W+�QŚӡ�ӷ��J
�M����%�t�0㉈�}�4ͨ!"�]�J"��޲�"�s~�GS��*�	b!Ds�UP5Y�0h�dz�HL��ZO�A���m��6�]X�O�ws��_ڃA�A�ឈ�V��ۂ0YY�fiH�(Lqu�i���7ON���sQDB;GĠ��N-I/F`U  Ǚ9��&��  D4����:TM1! :fMBH]�t`�TTRbdF��5��D�rO@ \�<d7���D6yt�b��[��j��2)Bb�Bf
�hvTU��ǶC��i�!��j������C�*b�tF�X��1%*�
�k|�m���f��.��0�-0(�@�c!ly�7���:5ts���g�K� �$
��|�&���
q��߾MP�E�zp��Xv��)# #i6!�O�?Õ��mK�@1�4P��p�!�Ĥۀ���0%I1�um$kD4hJ��~T3�M�m�tP�@o��WRJ�`Rb��Q��g��}Bp�s�e��WQժ����������F">9?y�����o�I���0U�+���/~�_���ݨ�&Dᚼ'ޤ��L�\AT��)���$hZ
⬵lRk���I ��&�'u>	39���<N�fFM��97��� c4V_a4E t����ܿ�j���3���~���O��f��d��;o���?o��c����O���/�.������?�gݺ�>���O?�Χ�NNN�����8�q�Z���/��?�aۅ�?��?��?�#c�`yC&��o���,���Y����  1 ]Q��N�T�y�S�1�cBª�-��y?�iYs@����c��8�U@"��ԋ�Ȣk\n�Z�	��0��ƞ�a��Rf�5�ڷ92*i�� �*�4�� �A-w] hSa���lho�+���8�J�R�A0;�H�dMF 1�Ϡ���Ĭ!c���۵MK�sj�����?������UB���l6���m[q�M&�����_�5>���nQ�={�e�IRBP$T�$� h88l|��3�Nm��L׶������
^�!Ѽ���\�|�$�me�H�YK6�$b�І�RmF�Y����P�!^3�عsxʭ�Ӻ[;�PE��<�u[#Y|J1%��"�mAA�V�fRk�i���P*�"��i]�܆��k�>�z�y�kv�
 �(����d�y����(D�H e�@U.J)�U1\^^>~����������l>_��$B�!�Rq2�1�c�'O�\..k_#QSW�C�}�d�'���Ն�� �@���m�r�B�E7�VO�Ĳ+|�c8�������6�XT%]{��o���,K��Ո�˟���)��esc��ҁ�;#3���7��G��̙`$6ڝEo���5�B�䤴	�!��x2��dBgk�-Ƕ4����TGR-*/W�i������c�(�Q�)�G(��R�l��ȷ�'�(��LLUU#*��ӱ�W@E��+_׎��XS�α�[�E!�d4�|")�"��v&2�l\�rg,�i��d襤yq�0F�������k�f�X�����콯|E��R�R|����{w}U=x����l<��/��'/�z��a�ZW�r�<�8�)M�#M҅��hI�b�H�䜍�r�4iݔ�l6��*	TbH������I�.�G��`⊠�Xa�4�9Jb.peb�d(Ң�\ٗ�!m�'�٧��3�e�Tb�뺪����x<v�<E�[��x��B��:�(����Ѹ�k�q��x�9l���tF��U��WU��f�Z��9��Ȇ�~b�)�+���s#��{�)���vx��1DM�f��/JťN�I �CaZ��Jn�7��,2�"f�1ի2%o�`V�=c�ZӪ�RSA��x2����y�A��kf�s�u�3�r�s
��cb�\]U����QPBbǚ�vIU�����t��R��5&��TY��-#�R,i%J�����WƼâ����1{Z���;-��9���%��3(kp���T C�CQ��RbO���@sT�y������ݙ�-P�$	�E�5��8�����VE��v�$)+Z�E��A�p���^��e�*��B"�T2b�����m�  ��4# ���OOO���9����'��x4I" B�������v�>���w&;/�?z�����yUW��$i�IL_o�%}El'Ԝ���sUIikVR�8��-OU"Q(A&av���n���*E
[j�C������(lV�nv���۾=��҉�v;���^�0��8��$Rv�$�e�`x�P����_<1^\�./ggg�I B��D̄���D0�,��;��ɧ��u5ݙ.s].�m��C�������z�Ͳ����ׁ����0����@v�2
�5/j���@o���xIB��w]g�����qJ�;���W׍	���'�MR��ԍ��ǄJJ���7sv�_ ����Ř��[.����{����!����!�*=���k�L�uMӄ����ݻg�5��Tк�L[��.//�8M��q3����)ģ���^����+����TS��,18"�5q��_,#�5T%���C�^Qr  �/�0���������pV�����b�*њ?���m����]��Jk:�
j�5I�Z�/..NNN>�䓳��:�z�J4) #����NOA�ijs��
�=��v�:b7n�� �W���?S�,b�c��N�5_��o��S<X��$�c�@ !d� ����
��HL9!֯z"1m�����挈��<��d�$wK�H*�6[��2ZUUׅh0[�T`Zu��J�B���-��|������ɓ㳳���Yq"C�&6�X9��NOOa9_,��3�P$��A�.�[�bq�a���a��KD�9��m2o�]�4X�IW��ˬ�Hk�KH4@
�1�x_ew�ܳ��)uo���\9��6��E);����qIb�uucMA��� ��]�1J�E�ΰk��1����ٳ����*C���43o��H�F�����"��_���~sE>�4�-� B�#oQ�޸V��DIRUUE-�?>����"!y�www��njI	PG�QUW���@��BJ2��?ΎE��ӧ6�f40�[;=���O��_��,R���U���F�Q66�K���f��7�K P�\*��DRLѡ#�R�� �b"ʱlL��@��WȹLXȈX�ô�;"m��w�me���Q�M�y�
D��JB���c�����V�hO�u3z�����s�ᣏ>���O�j����dg�`�1�,�����?{~r�eS�MӰ#fJ)��yя�d��&�]�`�]_��aH�yu�e���O؞���f�_6�Ԥ^!���Iz�,��u�g0�@fj��Li}e7"42	@
A�͙�0��5�l� �c"䀹��j�Z,����ժ�X�g��Dq��h42��/��1�Э�.��v{g9�.�>|�W>�����p�K���#!y�lp��#&H�˛����1n��/*F��m�Ŧ�������l�{[b���t(0h�G� ��� %
W%���'�gg!���ˋ�,�xpp����R�L�SEDٱ����������񗏿�G��_UUurrb��iwa+:�U*��k�m�0�o�q)����|���}�q�xK����n��4fe"$6tUTgD[ь��G�($�m�-y#;"�x�[�c���si���F%� b��"&���|��_Qq>�_\\ܿ�`wozpp`9
)E{`��3�z�^��Ϟ=;~�+TX�V���"Fus��&PN��Ѝ���I v�/CP�,��f���u�; �� ��V0ǟ28��!���Zm�F�%I��X���(��4�L�ꋜ`c��-*$��s����m����g�V���d�mP0R��^	�S�-B�7Z(�	=���&�$!Y�I�hy�m�Y�[6�z�AAM�>'���E ,�"�&-��j���K�C xv"
���T��6%!DY�֋������*�.��}g�J!b﫪��]�"��6[Ã}�rk�?��J��=2QV��M��͇3��D��!n+�Bڎ��1_3�01����nv�,7�?��Q�漢��Q-����\a��Σ%trK@@��9rP�f.	�+o���MM0�놷6t���U� 9����Ν;�hy���#P ��R��vDE������M�I�eï��֬�\�>{�r6�+.�/�h�D����Y+(�]����z�\.b�*��b1P�
�4)��q�1��n�X<7)���ds%����h4�@�1��M��N�� �aT�#1���h4�N��K)��z՚h(6uszr����GM���)��n}qq�� "���+$% �y���&��K�^����.�mGc��ϥ�������Z�Z���ʫ��Y��b�s %�y�4+�@D��/��������� 3�uSU�L�={��_�V��jyzzJD�y�<"�5l �1Q��(� �TM�j˾�?m���L�[&X�����+�5H�\��lo�$z���썧BvzUͼ�0n��_�[����E��X (P���?U)�k�r'D@�Z����ML�M^4�Գ�{�6;QJ��"Bg�����^z�d���
!��Y{ɺ���L��/�<y�u�z�
!�VK k��@��/s�H�Ըn��?d�X!�n��u����oxO�V�*QNR�h�EdE8�і�E��qQq�� I�<~ظ�6�{�D$6�d/W��u��3�}&�lp�&6fY���ID;vlͯ���
7a0 "��4d��s�����,-3��|�ྯ��j�/n��ЉA�)�e�I��6^p?p=���,3"���5�7ճS��r��8/&�~f&k�q�`hC��y7��+���+ɘ�aZ����l�PZ���C`���*���#��p.CQU�\�P�Y�7�L���h���� Hλ���V�.;�&)0��~M�Ӡ�PVts9�ݥ+��-�W����	�[�6ل摈(1gy6����b�}EL1B*�c
]�Vu
V��"�Vh�FV�l�c����2���t�~��i���)#�`o�5Bo
��=}�ѿ+��  �(7_�L��,�h�~�QE�*� X�=��$&M,׫��<�X:���� ��픙'��d2�1�mk~a���J^,BNZ�4�º��jGD���/^����aU�"0xv'�'�G�G��1%f�kc$U��_6�،��9̃�A(��C�W�Yos�f�?ݏ�kRh���7<�fee|(/����U3�:�roCY��������3�H���m�wEk�� �.$��:�ѭMq�3��i;H�Fs10.C��Ĝ^{�Xb��}���E�۬;�/�ńmTI��g�� !211%�9�i�r8D���f%Sb�b�@-�`��#r�.JT���e���b�����旼��T�	�v7cE�?��*RaO��Y��U�����j��ٳ���:�낪�EbUWL$���zvyم�0����2��ثB.*�A�8�v�@4w��u�u]��Ě!�n{	�D����V&?�U��[xS���>Iz�M/�,Q?�)�r�-��(��I����GR!���MSWU�-[�� ?!!
9竪a�1Y�Ҽ������"���B��9.��X̲o ɍE"D�XM���x�A���~��RC����w17�̟�҇ ����a�^4�إ�%��FL"����$_�ۯn��`9�!��aB�\����ev���:_U�����-cU�{�ܸ�n�4e.�->��Ɍ����y�,T��}џ�`����x��-s�Ϩ�9��DZ���n����*̸`��s̅ggg''1&(�^��mN)8��o\�d: %��oH2��ޛ�F�׷g� s.���v�����O	�7VfS6,���x�>w���yy؅�-7`"U��� o[�*Bn���qSը�!�FeAR$H�4��dǮx�Wc�|7���E'��xn��12�X���5t�a��7oT�B�������`ww�i��3�B罳b��RL1t�l1!�f��X���-ϸ�&�'����dt���o����<ѡS��ݙ�vA�u�W}����W��p�nj�z�=�LK��P0�b8;;].����D"P�QT��M۶3	�<v���*)��5���N7���p��v������i� pq�t��Ӏ3L1夶Ew�������à�\¥�w��M� INfn�\%�L�`�q�$)w��FT�������̌
�DD % u�p��*xgIeq�mlW����1����s)@t�!�*"��cN�, (��6 ��}�<u7J��^�*e;͟)+������X
���Ke���VU #�O�P��	��J�=��h������RX"���Ŝ�v.g� jV�GU@TA!dU@r1���&�Ȉ4�ZG��,\��/�(UM�,�C�d��n� �)�yY�Oz�U9o�xuU��l`���}q�O�������'����8E$1K���s�z1U��1'*�C������1X?
�T����>���j/�T�@�����Z��z�@���J�-�dm�?&��R��k/�Ü�0�G٘6��j��K�k�������FTT$���20;��"R�v��򻺤��%x��+bp��9�)����|睊&Q)}��Y��Rޛ�0��>����kK�b��=�H��WQD�2'I�
.6k.����Z��تŹ���H�"Iz*�#Όgn
��?�hҤ�}�!���5+ԣZ" �Y?S��MW ��I��~#U�CYݼ�,�mIR���*�8�zC	/���y�Y�g�e�u��zwwz�޽gώ�l�uU�1SS7M�TU�*1��;GV������pS�����8�������_�@t�U2t+�WT���p�v�=�vn1-��� �c����@	TՄ�c��NN4��-vs�%��A���ƕ�l>�'�o+��Ԑۺ��zh��  `侱9rQ����7��(fe���R��E�DA9gz	��m�x_a�H�ڃz�����r�� �66�hm��LU8K1Z�1JT�(d��/*)R��;CpDA��+}� [GDE�NR�&Q�5%̲
�`0�Фػ���Oh��IELTu3�u\So��7$' �K@�{��-݂����%-��H�t�t�t���}����|�{������Q�5�)j�ҭ��4��ntl�S���_�I��5���Z�ǋ���?�~@�"/�"	  ej\3�4��ڎ˞AXl����_0!vj��>0�\IK�c6dIki`�I!�M���fƏh�;
�9ߑ���B}��7����w,-v�U���[�v�Y;�M�@���Tǘ�/LΘx`j��Y0Lt'�-
��fOX�&�m�?��t�?�k��C���Y��E��f�B�ؕ}bp>�?�l|�Z�5&�䦀�z�U�c�8�$����89�+�����L�_g�>�j��ܻ/'��QI�1�������pw��y�h�� ?+��I&U�(���D�FIW_V7D۵r7���4���~���5,�zл�{�`�o~8�kΉ���O�k��d�$m���Z��uN�Q�`��0aZ�J���	�K�6���	&�4�f�P΀g��ux-_�V�B,�����ß�x��O	��L���OM��y%�?��r����t�"Y���1 N������
�n������ٲp�>�44���`��������qJ�u��&�M$�
�c�vu�*�6B%��4��5U���|�G�ʑ��_����(&Z�Rlk���}�3v�H��Y׾�^�l7ҳP�"$j�L�ӳL�k�<�#3����}IC�3�d���|����E����x����+�[��W˱>�-Hm5F�8�J�N��Ў��~�F.�%$$/r(�U꿑�_��uE�M�d\����[���8���ZߴL��+j=H�AZ.o�T�yX]-���9J*�|�T�hX:�J�1Nlɜ��>w���/]nX��A@4����,3����s�c��u�̗>|z�'ީ�6D� �^�^e�M!ջfW�{PX��돣|�MĂ:�7�o�F~�(q���9���p\=ٿQ		�2�� ��UN45v)�(N���r�V�n3����'"��0˯1p:^9K�h����-���6�u?�E>׾���U�}�sݢ(zV�m�#�9�%h6��>��v����'l�Rhp��S�Ȥ��j�P�۾�k�BCV�!u����f_�j�@&���}�8_=�ӆ�[8��Q�,O��N]a%Mp�{�R.U��Z��57eϧ��{ھ�l��'���#�o��eM��m�-+��u*�..q����g-��vr��,�U��H8�����F��Hi�8+v�z��2���1m%D�ۦ�M�+֊��IX7��=�p��������	>c���������s��v���[~ ƶO���_4�ݞC�D>B�\h��g�2��k��J�RIu�R)��a0��W�e��<QZ��l_���o7$��tA����.a�g�^�z�wfoh|��MH
K�m�G:R&�9�h�P�W{��nG�A�%�1҉&�� ��v��������Qq��_���S	���05�%�?�{a٩��;,��Wh�%΍&�֟a�]s>�/~��+���R�I�=����du��}I�Xwf�[�6�o�WKM�3�֣��?�o��
�-�h|�2v�.�]�{�Č�d��klv٣��N0&��������X����g�����}��8��a4WH	m��nL�y��1l��X�B�?X�q<0�����(K���I3�TH���K�]���Z����S�vf�QƣB�ZQ���XI݂#�@�Qv�,�RUG�z�1�t�n�&��M���t�3�5`,��5�/L�}�8�|� �Ge:2��:�w��r��w]W�\ԇ�{tw��!$���?�����F�Q��ec��� ���puT�����fvz�|;'�O-�y~0�ǲDq��Z��7G�Lӓݖl�N�48	��J�X-)�s�� (@�F��9i3�[9E�D�ǲ�N�8�AG�!��.�lϡ�?���	�kP�{N�Hf�y<!�z%P*���rO�%^�k!A�E~�MD���[�1���/.!!�+r�p�i֥��<����?p��NS+P�Ag��a�1�R򪜴IV�b�|�����{5��n�`�Ms�������y� �b�-�WJufꯌ���s$�ˤ�*�Z����N�gʀ��w>W�Z����w�:
ν�|����4w%�k�_�T,Ń��7�5��a��S�mJ"Q���55X�F�D�/T"��6_��
�)�8�2��[3��:Я�ɬ�-Tc�uV��A.Q������9 �r2��
�_�98��v�َcTâ@�W�Y2C�0+�,��%6\���kK�X���Q�U;,v���z\��&�-�WTqL��-�,��׌)P�����bv6��Y��`)�=K^^��Dc��R��TJ�+���4���֕�|�/�29���\��q��+X��f���}c�l�tԳ�ː���7�*y�N�R�c���{����ע��/'� �D(Jb�9���R�]p�	�A\C&�[]�W{�蒖�WWW�ְB��t'���kCM]]��_F������;�V����^�2�Q��%@�:�C	���&�M��ַ��L��+^�̎aV�f&�O��΅deā�7z����ӚT��g�6������l�&>6x�x4��T�19ῳ�h�,��QuN�����W���19|�����h
���"jSk8�����RO�'|��<+a��`s`BdE���9|�IQ5.~0�}2
uR(���@����0�ղG���ʫ�T~DR�����o[�?���H$JG�NU�]����0C�x���W�B3��Sf^XH���w�՟�ݾ�P��
�B:Z������;���Ff/�o�2c��ر1��<n�Z�s$�XC=~��o�n!�$�1
�~�O�,ugw��　�G�z�����F�8���7��:�΍����g<U�V̳�q�T�c',���n_���y�`;߫R")1�Wh�K���p���ǐcot���t´,93���U��Eg�Nc���zrii颳��/C�+dg�mD'��Iz��j�<�*�p+4�Xn�I:���,C�f:k۠��Qr��"'-�.w6AG���	35*�_�o��Q��T�wY6&�U)X�?�ݥ�;d�Kн@,������x���l�/A�l��>� 2g�JO�?���c�.��X���{o�;.���)���l��ϣɢY����K��
w߫ˣ�γ�����+�7�3F���tIER�.zogN3n� �>Z`�4���X����O(��M��=t0F���A�Ԏ��M��U����SZ�t3}3���-�T6�/��x��i
L26���>�W��[V�,��~�?ò�{�k�jY�R�'�� �}$�:�;Ml3�H>���m�3ť��"�d�ޫG�m�;��ѿ�;]kҦ��q��n%�wwwW~"���{ff����!j���J�6-���c&���^���i�s����2��|��RB?`��髲�ɷ��rGf��$����'�w�ƇQ.���R�gN�Eer������^ee`�㣼~�F�T	��<���f#YE���b�s1(Igf��=_N�U�OsKv4�|�֖c���h�H���S0)�YS�r5:��E:��eF��� ��SyD-nz�Q��3gnY�p�����>��?��us���W;-/,1}X�b���|%�."����1���g9����@'���x�����pM
��Եup��XA�ںA-�N��A���RzK��+�)�����{3�!�H�Wj>�d Y��D�o@��A���'��<;�`̿ /���[lE-9D��JT��a�dLE��ڵ1`�zY�F�%3U'4�$B��s��Gvt�%[wwwn��Ͻap66���l^+tĶ��뾢��+�I�&�����[G�����	�����ۓ߭��V��F���\Rt,�Z��=�!ֶ��C�t�nM�@�N��{���b���b�E�� ��1۲?[=?�׎����|�0�t1M]Ee~Z>Rۉ���9+w���	�Z��WM�h�������Q�W���Y�(0�C ��#��=�t?�E��g������>&D3O�昭]�R(t;�:�@gܶPK�Ǌ5 h0)���t^juuu�+��֗�k��6'O��狜f�����Z�w$���K�(���������ޫ��r�D�U���
	+x?�i�^�����k1����f�Xw0@L��g�ш��[�O�J$g��J��ߙ�ߑI�2��;]ږ���n^�S��?�Iv0Py'oP#嗍Y��B;�qn�ejdHx��3��ˏh-�Ը���F���C��Ɨp�����?5���7m��ss]W3{�.�O�ɍׅdC�������#p=%��[yp������O�i҅�xù���i�b\���_�=}	�B��0�#y���(�ӎ�����:��Q�P��v�v��8b�my_��:�m�}!�Z7�N��:�����.Z�"�����X�Ǐ�'/�|����ԭ%@mx�١2����;���I�x�2'z��"bX,�6�����׍�%���Y�����i8�䎖�R��g9��F�~Fi۞��v��H��x�0p|B�4�����͈���>�Z:�8�1�S.����-�D/E�9ȑFhm�up����M�^��@{S�� l}P��K]^������$:�@�,"�g[��h�P�̶H�[è)-!���W�(�Liy{_?���s�
�7�'!)*�W�[Z�����#��]
%�n�oՐ�j)a���rua�����o#�(1)��8�ǐS�v����{��=�r|Ha�τ�a%%-êH�6W2e�����\d_9�l=|�����F��<kצ�z'���y0�Gr��O�D�RN?�E��]��H*䱫�	���ꢔs["��+�)��R�%c��d�Ρ�Yͼ}3��YQtL	՚y'2���ށ:@}�UC��#gX�S^��X ' [����>�Ѷi�Clm���AA3�����hi�A�Z�uu���C��̐�6_�(e,ʟ�� =sSS�y�/+�P�$�8���Ko �Y- ͈H_�4��Iz��A�c���z|���y�g��`|<�QG\�0Y��j�C�Fc�C������ut�y�vT��w{���k�'�4m��&�F�Ͻ�2�z��`�� ^z��\�֘�eד���2Zm���^+�)lt8���#_|f���5ލ��k߬����~Ѣ��$��s�xU1�7p^�b���B����6-z	5Fݐa���VR�u7==z�:��:N����\o}����׋�t�dP������Z_�VqD�Fn��L�?�zt| �$�jģ�X��� ���Y ��m�$2�"kx=��'[���;4C��r;4�?d'D+p� >�r�P���Iv���8��f��p+�TK��v_�I6�B�뿟G�|iu��H���6���V��U2bs�4��4����!&죱�HU�"���a�B����ў<� y� j>�X:}3 ?é���][�
�%k��d4�:ІY�{��,	<�]]]%%%���0��zx��0XK=O�ڀ�EIZ��� S5z쯿]������7t�f�6�L�����{l��$F��P:�9�7��RܝSᖭ8�fn!L]\*�*V�9��e�������śő���ġߔ���P�������x��u�]s�2(��c�z����c�t�����Ntt����l���j�<o�j$��)�Ez0X����)�*<���>�6�P%��͐��A�[� غ��A[m��Փ��<UGoZS��;�}ʒ����z�y�D�[����X\ny7�� `T�-
�k�OଵƱsol�1���ՎG�Es{Q��;;�$�X!��yn'�I��'��˶����]#��GEM(��6��U2�"���wC+�����ݾ}�}����ߍ��<�:�+�����v����V�VT�6r2N��aT��2� j�V����#Eo��
|Mė����9�}���&&'���l�sTYf&z*o.׍'��!��^��F��B�|���BA)��)a�N��
�`����R��:F���}U��[�`A�:�zf�k�40�@��[.�F�.�,����aR�N!:Z>/����W8�Ӵx��i-@MKG���.T��U����>s�����4��h���lf���`^��Ձ����� ������2Q�����/e�ڸƮ �$YSw���y�`~���wμfұr-#�b�$.�3S"'t��G�	u�յ��?�nf���އE�op�VH�J��讀	S��HT�)����`�fo��)O��l��z����-�9��+p�b�<�`#g���[�%�R!#�%��'���U���Á�'~��6�-.N-Ev/_���BB�LMM�l��P(Tl�\��uy.p2��s+/4�T]������w~^�|&����՟���y�e�������u]cq1Tq�f?eic��bf�~������H��j�Y�MU��am��3�ЄzEw���#默yD���@Ͽ�%��ڛۄv�%��3�.��S,�8a�q�WQ��3X�7�<���dK1�% ����a賧�7Y��nO�J�^bt��l���\�{�D��	^A�v���~�JA$������j�"Q��,�ٖ�]a�J!�@e4R�bx�|=��1$A6�;A'm"Y1�a�̄�\��3�������1%@�"2v��K���3��n��"�� *֢+��z}���ͯ[�h-ǃ������� �803������ޟ�2�$���V�5�٪���^{�kJ�� &���6ZE��+	�t�:���x���~r���Z�.`�뜝�5��x�Y��3���� �!������7�d������WN�c��$�ꭝ]`�}n�S�ƫj����`�k��,����5�Nx��վ��C��]������Q٭��g=�ɮ��!�v]o�9SQKͳ���<��b��*�E������Ɉ��[��c�׆� �W�\r�H)�&+j�Yt>�����3gwRb����S�<9I�y%�˰39�Q$���dLT�*P(�2k�O���m���I3^P}KX�T�$�;�l-�i�2$6R��=&�R�6�BL�Qc �5!J���	,�A�Uց���~�;%)T��d��v?ʗ����9��X��fD�,,O��)Hƃ�E����-||�Rd"I��Sq�z�A��YVo��`�N�Oq�C�&"w`�s5gLY�-�1��X����D�S�F�	�ϛw�lQ�Su��~��"TP������UѸ������>���޵��+:��!!�ե���\<�rB$u�ށ""$,����_^Y�(zxL��,|�Ժ���v��Uw���TayЫg~$&{&�/���o��9�@
�w^3<��y�D7���po��K�mW��D�:�ר���ɜ�}6�3�î�Q�}O|�e�PÁ���G���*W�����VW;��q���+�wkSF��HW+�Zzz&��g�՝v�0�8w䬀���� �WA秳��
�^0J]�qr:ؽ���6PZT�p���������x v�- }��x�	��eӦ�f�Q6���r^�E4wq��WjJ�F@�,��J�O��ˬ���$к�f��5�azFK=9%&:��E[�b�M�ͥM��	2[na�����0�x����(1[��U2�/�
�ӑ�`q��H���p/��)��o'���*x�~g��1=������?��@�MY��\_�nn}}n�B �t�@�G�Ł�)���Q/1���P;�L���{SX���Z�K't�4Z�
V�)��f��w�m<�Y��I�="��;�u}�SI�"�'����Uġ���!:�e�OQ5Ѫ�F��&~��{n�3�w�����20���]Kl^�)ŗ�K�_�S�K��읝��݊e�h������K�8�ƨ0��h�Rk-YZ�gڈ�XA.���'L��IJ�^��F	�	�L�LLL��<�A���TPPT�N�M-!�W�.��� �X����J
�.�(2|�=#��
B�����+�m��c�@ -�j`zcg���;F�k",L�1	����z�JD�OWG�J���0H�1(�ե����(��p�`�@��.�̫������g&���y}�,�NS������+o�r�8}�s}������$�nE!!�D���V/�)��$�aJ?���>�e��@�Η�u��8�H��y����Q|���wm9P~s��*I��x�n3�(��dH|Y<�L8������Ͼ=�˧�~�g�z�qz�>�!�lI�GC~��^R�-���QNE�Mj�Aq��c��9!��Z�vk��>��b�|�����<�5��FB�� ��K%�)��̳�g�n�	C��5�I����|��ś<�A��W��!;k��ƎV!ꄷ{����NЈ�r�9������
��K���w��;CPPWC�����ΤywPY{����Ηp���Z.��˽����'�ڼ���/v��'��r�KOF����^�y�t����a֗2��/�I��u����F�3N��q_G��L�$cD,0��0�T���`oo�n,[���S3�l��(�^�� 8#��� ֗�D��?\I�� ��$�<s)*��A�x���Ś�ܒ��&�W|:s��`e�X��'��zM\L[����S��RD�#�7V!(�XX+�6�Gi��ʾ!�F���[S�Z#��

���: {�6mvvU���ng]��a�EJL���,���)8�j�`���6��������^0N!�f� ��	��s�=�Vח��I��-����rR7vLQ���{�c*ց11����� R�Dbu߯���&A{z�9V\�U��z�=wW���C�MMDD��7���%Ђȴ�|����9��{�VHe���Gٴ��W�D,.�v($x3���}Wpw��~$�����\ }׿�e�������,l�C� 0*��jNQ7Fa$�7v׳�>���/9�ݞ��[�C4,�-u�^���#�9%
4��*���ۏ�B�濰U��P�j����+�$��y�G��H��Ds���5�UP &����^��#+�`�\kB%�\���l�O�%~b��h�� ����}�c��;�$��.9p�,lK�
�n�4��כ��;�P���e��)�L���$�������SY�+�T�u�J�Ћi�Ng� ���?��=C �S�433�=�(Όzf��5H[���_��]��M��P�����������Y����>�BB��D/98�Z���~֛uS%Ó���m��ƕN�lϞ:�e�2��PPP�^�+�+c�J:d��*m�X�.�w�!�EH�s�ǪU�I�i�Ë��9�u�Us��P�F��@�>%�d����~W='����U��o��ԁ2[�}�DQT���B��Z��DD'�+��-�a.�muɳo�kR�L���KQ�z����z�&ğҐmS_x_�Qny��ߊǽ�J���kkj �;�ւ�=\���=��ch��3�V�%n ����J/5�w��C�zZ�#��5Y$喫 `�o^S�Xz��P���"U5�Y���[���|�$w	��,�m��Ș�q���$�]��������y"⧩��i���0��"X�m*Ul�Y}���Z��!yu��10�0Ye�g� ���=nG�Ռ�\�A8ߴÕ��?��`��i
�O>c&O�E���Ŭa@(!eh�C����R�Ӫ�����^Ӹ����i7k���bC��vn��ւn/����R�_��}�.bk|�kiT�>��c} $�w:.<�h��L���(���~�|����w;�E�!!�Nw�����=�Gn�M��kC%��uIS�!�M�\���֩.�;���I4[�?���3ߐ�#���2;#�9�OԊ�|���fWcR��V�Z�Rٽ�?H����4)wg펋��g����%z{-�8���>Ȫ�# U�~��[LgL���OLp?���<�"�!JvM��ಶ���6�>�bs$U��*�\���Z`f*Q4�'��VF ��,'�dP�׻Ƹ��|!1�����K�@��|+�)����#���H�Xmص�`����;�^����b,_��0�SZ]8�:&ؐ�a�A�#��jrKZ_��t�޴�48�r:	č������;������HQX��ù�)��\�U^�IU��,�j�wr�
S=��P9v��t��̈́�9�D8E_P��l��+�gn�;�JĒ�����`$`Z���r�|+��� �������NQ��7o�9�n�n��t]�h���ni�
�

�>�iuX��)8:�5�7��_�������5���h�����$N�s�ԜԡJ+K^��r@Wz>��2YP���<d�?���Bh#GeM��q��qI�6D�ϑ�����۽��PVڅ�ɱ�F'��X��J66��p��$�L �Z�N���{���2u�RoہjVj��:d �fx��X^�����܍�k�*���?(kC��Uҧ"m�9'&'A{���.&�H{O++��7^^�q�����˴�l���|[[��:����I\����&�u��Wz�}:zZG	/�愅\�%�/ϛ&%�D%8+�	�~C�����o?����6�`w�dE�v�4�T�N��Vu�O�	i��ɶ���3ߝ~��ж�B�:�15�o�t�!7
�Z���hll��'C�
^�Ì����q����o� meZPM��.%*d���hZ6;Ɣ*�V���ύ�c-�sbyK写MD�����U6O�q��>r���%2�����0��lg�J�J2=�(o�p�Y�Fl}#�~�dkfn~�����T*uvuը�9���hԙ/�kl�>s�vћϨ� �*���Ɲ-O�Z���[g� �@VܸB};�l�͆�<Y7J8��4GG����^%2~Χ�>�K��5!ܝ�	�Xdm���\�y����V�	��7�d��Қ�����a����V�j����#�]�P5&3�~.'X4i``��L�����2}�H���OAr�_.��N��E�z�2�RSC#����Z`GA��R}��{���m	��-_ \���Ľf�}�ٵs��t �d2z��Dl���5g����"Ͳ���m*6����O���̞�{�e�E�����P�ӭ�(+J% #Ƌ�t{�ʹ$$�x'ֺK�U���2UX3n T�Y�AZ�Kt!g}�A���G[����M��-�~����݅�L['��8��Ey}8�h��vR����Ѳ�����N���Ŧ��p��Ӭ��j

���Z	����[�L��m�Y�<4�x
f�=��GK���M�����g[n�����z��|���'�^�ղv9+�~Ac&�k�,I���Ph�6�������u]��rr�*5���������Na�W��ێ���� �e:c����������T�G&��K�bJ2�����CP`p�U6��﫚�����`^��D'i%��J���/����o�����諒�7��
�K�R�Kİ���I���4~|F&q{�=���?���O�ؤ͍k���L�P�6u�S%=!�y��Ȃ.�#7������?�J��&�*p4��|I����l[b8JUc�a���;�9�io�F��1��XT��=|�`��Z�gUϾxe�����}�\�9N�u��k��/�P�����6����VX-�+B��Nr���B���>�g���,I�z\;�V]�9���*�Mo�T�$.�Q�����Z�y�=�	�ڧ�E��Cpn]VY�BO6����������Ɩ�hH����������������3�]BuGj����������"��q�$�W��[A~��''?]�XP?`�(�<#������L4�?���u��3#�k��{���ڬV$���X���2HH�j�eXᇩ���L�4�oj�݆ГL�捥�]��w1l���os�˭M�c�j��Ρ���c�77�x�i� ��_�Bஇi��^�����299������x�/�l�������v�O1	� Y�/E�-::ZY�6�p�?��|z!e,g���ƫ}��X|
%��f������㩔g���_����*
j@���RM (�9��TVYt.�����;��3#����o����Y؈� ��)cR�/�xp�׊XQ�Vz1��"F�1T��%�N�=�QYCTY��&�V%�|y2���
��o�ס��w�'\4��)��_(��p!'8��	���W7�if�%o�￻��7VR�{�{����	p���c���x��K�'&4�[�O�y�֤��@��`�IW[[�mB�f]S�����S>s��P�`޻"!����0���Û/��j��<3f�fi���V���C�:�o�Dp��܅�X�$wͬ�u&�*�j�mPc�]��pڥ���1�}������`x�@75��Lsa�w�Z%l�/��K�p��ؗFq_�_@�|����7��;��^�=�\��''#�bզ-�!���q�	��WBB,%o��̯�W�cIː����W�*=�	�Z��a#f��%D o�+tvq5�C��P\iX��Q̽o�ϙ�.۝�0�E��g���������j�F��խ^�;#C�d@:��q��Xj]��Q�ts��݄��%ק�d&ڹ��q��&�|ާ8`�Um�=0������:w��p�ߩKg��C8W0K�9Xʋ4��|�7|��9$�{!g֡֗��EԜ�do���6�<��e�$�y&;;O
HOG;��dip��LKK�QA!����P:�D�sss��|�]��Ӂg/�==�����
&�n�;�lg��P%���/���GH�A㋧�9S�t��a�.�>p��F{\���݊�C�������$Ω�ʈ1�l��Ӄl�E!4�I��+�ڈw$N+�Q~<M]VaB��7X�b�lM��9�V��H��Z�'�f���,ғmv&��Áz�;6�K��b�!��s�xww�&�����wS�>ů��D$E�P�|�k/~-m�D2��6��SW�c���X[��5_u�z����6�W	�R2*0��;Ћ�>�.�<���t0��y=y^}�ز���b��j�4
��幡,"��AL��.߉��$��t��lID�'َlQ�k��c�hCL2H�ٷ��}��
���o/V�I[��~f2�}���3"���:�̂��R<_�R�{H)���c(~��6�ٱ������o��qTT�@|2]����C���'�K~��Q`�V`'c7��-�s���=��a���_ѵ�j�G$�Xf�����+�TT�n�Ef���V�qk������Ǖ���\3[˞J6y^A��Ar�wk����]��7�YƂTGb%�&���1vh ��A�bX��!��tI�8H=L�E��uz�G�� �:̟���'�1ag���=9�������D����8c,r�6��ǬgmYJRLLB�~��mCw������Aϕ�F�K������--�U)����x<f]���"��V�����Y��!]�k�����',�#���g�p���^�^$�q%�|��S��Xs� &t��!���ǟUQr��ʐ��A 2~���������B���qy�p�s7*����	G�����(>�Vf*=�:�Dd��hJ�a��5}:���eOBn���).a�2�C�3O�o�k�t]Dw���|1��:��֪W�j��lx�!MﺨƏ�/�V�%r�y��	(X�Ώ6u0�~RJ$E��"d��&����{��)���)X:�w<n�_u֙�M�	�..�a��WcA~�����Ԡ��K���������p��i��ɔ`�ۢG�o�u�1,s����JF�(��؆�6��{R%f��Y%�9�-��4�E����K�2�Ր�? Y�3�M|�h���M*�� �`;�@�<Z�F�T�~fm�, ���H�OGǄ��Q���WBm��^E�ݎa�-O�wpp0�w��ׯŶ�� �����f���ȫ�@Ä���{#�F�>k�u.O���T��~��{�R._�������)��_.�=5���z�v�I�qb>�Qr4̃��Ub�ڰ��{Hm̘.��ݘ0;���1�-�gƩ�,��6ES|K�4q� ��Ex�l:+JF�3QT�fH:�W�K���4q��o^E�-�v��D_��Y}C$����~������`I�B>�*�M{���h
������=.�	�� F�����)*((c5��z�e�u-y�Z�=i}���Sm,�ml�n�����loo?=!�0#�#  Z]�+������-�r}e�?�(�.hA�eax ��^�7}���{�o��1<C˔KԢ�a��&��@v�GJK�b�yM���^c�G]|����sڈ��F� V�d���k7��x���q�D�i�k�!�?�.g�H�F�s���� �.���W��Q��a�ABn˗���76"D�����Q޸�x[[g]-�T^��ۛ�'P}�avv�+�K<�D3p�އK*��q�w�{���駊�x�3�oP$JA�L���=�힯�O*��\D=���k���+��¼@����ǘ �Mu�����4����-X��@tD�|/3;d��J��%ky}��__�JK�?���PSW�W��C�tcv�wH@C5����dw_��c:v����7\*��y���e�H
$ɴ�7�N�)�ے��|�����#��i�ה��M��ĿN+8��,�7�|sX��� �5~`����ь��P
��f���[��ڄ����/]��.�v�v&�Q(T@s�XѤ,p�bG���E�P���;4�ab;�r�;808�ę�i����B������L]_�'�lgb���*��Hm2�a�`|�^�>���#(��S즒Z�^.���E�����[�0j0�	�D�r�֒�O�Wo�M@�E�C&���SE�?H������2C�|(π���RG7[���ˊ��R��1ƈ������S�T	�&&y�C�p�N�P�4�-�P��K2U�s �](��`X�c��F��X������J�PO�X5�ߩABf=��y[��R%~s ������d�A��O�_�Y�)6����aej�I��R@1�^�o�;O� @㋹<�C~��
 $�*��8�HY3	3e)�i�)Z�u��7���?9Ɖ�?щ���*�/l�UZ�`a0�:-������"r�=�0�]'�џeB�EA`��Y��`���.�˽�pq�IR(�IK����ep9N�w3���#G�L �5������a~N��E-�K�k(����a�%����$�&lqV����%H���k�k�)�S��<C�Gy5�J�H��
���d�iY�J+	*���y�^��3�3���Q�aC)���s�0jS�Y�q�!g������u]:����������HJ���t�~'����5_��[]��
_�N�E�}Ss�����w�)�W�+��@�F�oe�#w��jQbTO��f���u�١!W~�0i��L���\Q;�@��H�^y4��U��a9�q&�;d�[�K�#Þ?�S1�,��,��ń�f�DF	PPB3?\$�fƐ�c���2GX�u����~=�aя��r�m����]�=�.8��cl9��W�>
E�9*R4�2r�"����7`�g�����Ϟ`g�u<C��E�>ľϹ�C�-��7�'w_z"|7���eEp��lh�\ ��߱biJ9j���!��@�f��^��Oy����i��Y{,����}��x��B�涺�����xm�r���;�����Y���uV}F�"n�Z�����1O~�!୏���|�)�wHim����3s�2'�}y5>c�p�����
f�O�bBy}^]%cX"��9ږ�3Cc ����� t�쒛���1�[��#�te�-���r��u�-�*���Y��1'O�~�ԣ�(�'�,�����|y_��M	�Md;�m)�'���R�!A;;�2V{̢�����t�rrxxX���+<�kw��x������=xim�4�޷�\tO~/m����ߟ����N%�@P�������9�؏���0��#�+�&�^@�hʻ��lt�?�B��N�d����8>1]���|�;¶�͘��,>��G�4q����3e�߆M������9ZV�~P�ynvWE*1z�H*��w۶�� �2Z�U�+�'�t�%X�����ͮ�{!�²?H��v�ʩ/��6�P��lR�P5�z6K�#�ť����)=��9Q��j�YQ0�}f��1$�9�,.��@��������7�{����Y4����gVq|~~~v~ޅ�3�q�<�w��Kq���p2�Aa�ؐȓs��Q~��
�S��O���jv��BH\k!����5�}�4�����.�ӯ�u[v�[�c��R����Ng��9����x�WT  ����&(h۶mۖ�]svq�g҈�[�!D$��n����o��޹.��OO-�\U�4���GE�!�c���S"�ꊝ�m�\�gcR�J�y.~�"f��.G@�R��k65��y�͚��h �z{�Z�� ��fq�)�\��s��*��Sط T5t��'���I>�f#$��"6y)����bK7O�D�scV�=�Pq\��ܾ#A^�x5�@1v�Wޯn�ll쬭LƓ���*!�G#;�_��~upttzz~>=g晴___�޻���银�K�D()�`ڣ^7Y	��(9z�l�yZʣ��L�^D���M���5"�9אָ�(��r��fӬ��XT��B#� @��x��@Dٱ�>�B�M�x���tj].�f�43NV&��8����˧Ϟ���a����b]�F���z3��{����ع�zT�����Z�_I#á.9��v
e�ԡ�����=�RنH��9ˎ���f���Z�* 	����l ��j�1-�A��py�kb��l�[��b-h�ʔ���7e"K���Q��x(�Į��l�21��m��ib��M��5W?��jZף����2;,P�*BZTDXP*�D!DW�]ם�|��g!ƮkE�������q]����˗{{{�++U�1:@�"�SWdY�)�.a!��c2ȉ ��
"3�䥔�4'�0����{EA��M׵�P�����
uH�ET�"�]D$�s� F��Ƅ��$d$�h��dE&��ʮS2�Z)��2;k��L[u�$�͖�B/H:"Q�k"��b���.�F @4�K"$�,�]g2׈�Kkڶi��x���@w�����h�D�$bH� �̀Q�O���2Ac�O�����p?[��̳��X����{�lLu�ёU���T>"���G?�ڕ�.B�C(:�M���h1���|^����"�*���ATT@��k�|����:�kT]ɿ�)������"��޶���{7��1�Xu�)f&��e"[�0��ݙ�gK�y���7c5���E�ְFFb�(F��s��E4�I�����HL�9@p�9 ���h#�1A{;����;.M�Yڦ��t"�L��*�cu�;s�4�K��&1��Rc�$Z�g߹�|ш�8��r�@���H4��`���b��@F������g�J�̩���z]�������J�Dk�Ӷ��n���G+��Cf�=xw���˯��͗_�x�������~��������W/��2�@�@��k'`0�j�}�N*� �*�s�����خ�Z����"���9W,�c!0�R-�cv,*���!�(*�%_BS1�PB ���������[;;��l6;==�m_}���4m;������4���u1 �w����E� �2�H��[���} ���ڕy����}1{H*�s����Ų���2r����˼4��~���J//��D#������n�d�Z�s�,���1b��t�1;D�y�Jh�2��� ����xU��D�h2j8sDD�sޯ�L��7@�˯����D��l�X,T����tέ�����lnnp�0�o�1�����/'+��fqN�����`I�A�e)���K!�A��D��?#5ƈ��&�=�n 3v���*��ل�q`�w�⼋1��Vo�r9NE����u��(ifsb*�#$1�O��i�{M��-�UIA�R)�Y׬���R�{,����y�" �>�	�L�qͬ�QD^��\��1t��0Y�:�y5S�Ĕ���v�[,A���Ҷ7x���]{+� &��{�%�j����H5��(��\�c�)ab#@ȁ���E@�"��o�Z�hJ���ךg2 	س��*`%��l�����d�����R��_43��I�f,�;�n���hզf\�����􄅳5�-�V�J$�.rT�Q ����;U��(QDYS� hb Hc���sN�(Q�M}��ܧl��DB&���WEQ�� � �%D�aZ*Bz��H�a6:"��$6\d�D^�6p
&$0�x?0�����%g\k]jQ�Ҳ#���2 #�j��ҫ�N�2�s�y�5b/K��wo���19"E۶���f�3;�{N�OH�~��?��W�*tag{������hc}�޽w��" �կu|zrxp�%���;;����E�g*2&W����q���^!!DQk$���'E��� �YtP@@&R�����  �`Y\���e{rr3��J�	��!�FTt�����왣F�L�J������/���s��k����ߏ! �hd�B��"9W�tms�s\U��޲��:��N�[-�č5�>\�r��I���j<�!��4a�CQ�K�KNڛ3i���$@���5�)��)K��Bd��� -q�R�$3��[d4W
�b�T'b@M-pz�	{xHP  3�Y		�X��1�&%vw����?��ի�UUUU}vvv�Ν�l�������}�ݝ�[_|���d2�)�.�;-�V:dY��JX���>Nޙ�*1��j�6��T��͝#�.��Ѐ�0�7ex��&�(�~DpL��s� 1�.�m��.��-��*M��p�$�u)I!/:@˿�!2;��J)T�ToI��r���h	fV�� H�
���R2�!F����^ ���E_�۲b3�
����F���}U1��s���)+�I��)c�]�l�\C���9F��aO��vş[>,�o_U���-uB@�V�l]>���q�뤑(#V0����D.��i	",/EH����ù�)��{�-��	\GB��0'�-Ðf�8z���
����CQ'Q��C�R[t��{NXR���s���Ѩm�Fs�bF��!)�5�'��J���)
!&��eLL��?͖�iT*5�RJ�A5����i�T��c����4�50�f2����ܨ�G��������>s�_:k�HaM�{�-��#��J� �b*��|�AB@f6�f/�Xa��� 	��Yĥ�r�ԡNu�!��� ]�P9vLl�59o�{!�Pޫ�8�DV��HA����!!:գŬi����۷n���/�����sG��]h�ݻ� �o��u������������O�O�O����.t�H���Ê�w�Q�^��|�K�)`�{e�u��8㉹�AT�}�E��2Є�� U!�+ET˚Eb�\�
��Dg�� "�KD
�CAUƓz<����	���h�w0X���\�i���s0��p���Y_��j�c���
�� ޫN�-��M��Wʌ&���b�dV���g�>����� �}xIW� A0b�\Lֲ��vD����W3�B�{{�
�HU�R� ��:Zʌ�CU��:��7O����έ��w�4ms��} 8;;����������h4���z�p���X��Q�̝�EkNQ�ג9\h4�F�#�M��] ��Yr��Җ����{��9'
�:,��U�0JT$�Q��sU]e�%�!�F�1�Hw^��s��@�Vm�~Vr�"RbD��U�F��8�r'D:b7,o%T�=ʭ	��s�.��W�]M(eN��D�H݉%�[c�jV۷D�l�\d��1�AqD�#�0J$�wVZو�"����*(���@BJ=#@�V�A�l'ke"�h(��q�b>$((�"�- UwE|) ����O4�	�ߦie�[ �BĪ� S:%# ��J��1w���:ּ��Q��+��Z(T�cv�jq������ʭ�(�@2G�1�.��X,��i�6������IE�� i#��C��6�Zrj�B��?��T�	Q�_��B*�<I���u����F{���1̉3����[+1�B�2�GR� ���a�?��H�� u�:ϑ��c��S\ZO�'�Ք�w-YUȴ��k���b P�C!��i��QcW!(�k���Bwڞ5mc=*C���|�A=�~��t�h\���E����?lll����;9>:?��LF�J�\�~�o��"J�Yo����99R����R(���ǈȎ�Ē5x�1,��0;��r�4��K!y k�ys廧G��
<tM{�A��-P�A�M��E!���RK���Y$R�pJ�<���^g:FUb��K�4����WC$B1�/�T1�� �e�AQ�^�-w�sQ�D����Ja��2�})d��|i�m�D0Ah��Y�I����V/��X2�ND2j�i��FQ����A?D]�j���}��u����V����������d<n�ֺˎꑨ�OVХ�)�A(�e��
QJ�Ť,�br�ȹ����7~$+N�^0� ���bᣵ���� Q�k���^At�Y#��� ���ʷ��\"�B�h�8C+�]^2e���2l3G��+���cB�3W�*�^l��4��{/�=���)��,t�����ὡ6�Ç �"��Č1v!,�E��1frv�Y�?k����%�ȱ%b
��8%�OD�=NjL�A4I��N>�y��]�ɂ��3��b�\�� D�z�o�Ra:H@'�� ��ypP��l�^�B@T��h� kW�2�B0J `��4�_\�R����s��$`nVd�J�zp���Oq�۶�M����EE4�(9>�*��"�EԠJ��KfG̈V��%K=	��̧z@��O)u�BB葭� f�,}���d�������6hDR�W�<��X/
�ۻSE��+�JDQ�\������7�|;\�N `DϬ!�"�\�X�5W6��&���I%��ta�a�ݷ7���[Q�WAH~����^���yn�X��b��u%""qss�ywq1���M��g��8�'�}����������KUM[= ����͓�;�,c�f��Hu��i�z�.k@D����l6�y�i���I.23���PPo�
~���������)�6���v�I�ر�{�������J��W~��iY� ��,  �ݖq�c��P�ԐX0 ��r�[�a��~K�8j��F�� oM�����������!�8Ġ��/ƨ"����� ��G"��|F�Ɏsb1�̢Je��A ^
�`��'"�g��=���"ĈM�vm;�WWV��v�ONOM��7c.JP��LK���E���,�6�z*�D���f<�A�K�& ���v�l6�2��6D�%:&�����tE*_%��Ɂ#b�B���@J䪪2�ci���]ׅA#�#v� ]�� ,b�X���1�YQ�U@)?��O�Â��G+3�����������<4�����h�A���Q)�Fa>�ϛ�w��.�	��D�[�Y_�����k���Z�1t!�^/��Sx�[^�~��O�^O�����Z6~B݉@R��j!�%��X�h.Х���\U�!�Y�;d�_�*�\6�.YƚCa���ָ����M9�;Z�Ů�P������VLa2��ΐ,V� �r��-'AɃ��2sN�&O�3��� 2ew^����_��"��C���V�V	�(���%zc��0g5�e��r�:�� ��~ڔv�`z�loq( Z�O�p�&�x�D��(�N,ex���e��8��Ŏ�P�J�N5�`Ap����\_���6��9캒Hj�qeu�.��b��+㕮�ڶedbn�f>_��{U��������ѻ�}��>��lzg����渞��'?}��y]�F�"*֤@�*Q�cY�>F�O ���-lO�N w.x-��s��ж���!2�JE�W��}�s�=�B����b6�4ヷ{�4Z�>s��k����|HD�߻1�J?�K��w]��䈚9W��(g��1��U�$_.��v�UeM��\� �C4�h0������*�@L��Vo�jE�;fHD	*"1h�|6�k罈P"�6�]�a��B�W{{����Y�s����b������	��G��Uϟ�8;;=?�x��>�J�!�`�&c��+6e��I)����3���*��a����:0\$�X�
�J�؅R�p)R����sH-@Bpu��0�/ܔb�U]�����|�,�:αs��+@�u]ۍ�瀅��؜wCh4�)Qk�l�)�D
"*	�q��ROL�����]0�v��c^��6�����9����+�X벁d�Ԙ �loj�	��OP�ՔEժDj2t�`u����_��u]W�`���{w�,��x�y�=���A���xYJ����V���G�?�������˪r��*H�߸�-���o
��8��[�/]	��&��d���A�;v:���lVG#}n��&���]����$���+�O��e!��)@j^z��^g	�ޞӬ�R�^�_�^Y�e��Y�Y�`���jLd=�����pxF1�B�kD�LњgcT	��JD�" TĢ*Q�Y�v��㰩�"QTUI̦��0AQUB�<;vH�_�j�o�?�~kϒo����hcXWս�w/�/>��sP]][;?;���C�uM�޹s��Ɠ��*��Ʀs���{w�5]AB���?������^��ELr���i�{ӛ�.Z{*FB�]�q"28�mZ�(�[ZDd�;�ED�[U�IT��QQ��9N5���-y/�ĵM+^]��}A�ܞ~d.>�!�!��e�� �!�������K��K�Y�t�Sz7~�>��Cg�o*�ϐ ���UU�I1�J7k�g^D2�1O�3w!��s�;g=f(5�1�4��iZ�X��NL���D��t�U�i���9�j������Ã�)*���AI�o�Ɯ��hB�1hnbU8LbREU�b�lذ�
F%E�PD���$�ʂ!�(F�����g�<mUar̡��vѴ��@��eb]�UU!�� �L�Fc?���5z��x���I�E�D/�L@��0�0�NA4���T|�VN�����&|慠��ĩ��v��P��޴�
�c1*�t��I�'���O�&U̩]�g+B������"r��"3S9�lP9��5:@ON St4���yD��v6��Ki��1eݛ�ߞ\D�*�$��H�(�LJL���,o�k��\��P#�dg���Ͽˡ)�nz�K�����}�b�&Գ\�&q�����y�� �C�Ĭ*]�%�`U�l���� �H�4���m[���C�r��/��&.�)�#Ũ,��R^Dz ��0����s@$��1�OG��YE���5�ƣ��5|�#��/��R(~K�\K�H����*Dg���"�u� ����Kқ�bNB@CR8�n�:OJ��29��ҢUEգc"��n��b� �Q�&�������[���U�Eۅ�|Q������b������4�ӧO�����㣕�h��Ν�;�|�I��ի��bC�LF�^�������Y��6���퇤�u�������sn>�kFD�{�%s4D��1 X)`�=����w?p)�x9Sd�j*��~�"�eeK�r�(CG8h��k����� &T$Mm�.�ZE���I�b�]�B��]�$0Q�X�V.Oj/���XV��&�H���4hј�и��'�"ڵ�I��!+x���TL1Z���
)F`��C�vF�}��F@�瀈��y
$��>@)���w�\�< @�Q�d�Pi�i��&d A!�j��x�"D��J�س1RA|j����.�#�C�C:D���� A��#��H�������NT�]A���U������%�mk4�h��&��x#�v�: �/վD�"6/3���3��!˕ĉ󚥘��BOuI	��E��̙�(�mCT��,�hV�ŋL3��H�����Y�hTS�!Ɣ�A�ȚڒJ!v�ų��͢�:�Ԛ�@�i
�ea�!��k)'���
&,n���-6V�d�b��׍f�qU�V2E�5��.�=������x��&f�f�c�$/�^��B���Y��%.�i�P 8�b��9�#[))
��x߈*�l0��땩I��LL��`��bZ��Vа#�	�N�T^S,�l�� \/�-  PJM�s�����('� E��o]=(= (-A8�&:���&9�C:�2Zf��;o��ݚ����S�"����f��@�[�W!�(^C�vcc��������^�|�������sQDWyD�[/������xTU�B8<<�����x���"PU���j=���޽{���0�൲�_z���7�����g��T k3MhhnBc,��oo$����Jig��x<�?d]C�&
$Qm�N�s¢iF������`�}��(��w��.�����8�`�䞕/R� �YaI����n8�@��].;|�f��W޻�5��g��!J�,=�s����qjbJڳ{�K�B�>{�ԁ�*�5!�*1ƶm�fѶ�p�iY ��Ц��cb!t�_�B�|�x�` !f �'��OK�9�E5/VH�$=� �0�b�����q�l˖I�\:"�;�����6�w��d4A6F�L�,[Z$�UU�"d���dX���̘,XUp]�v>�;��9�^9`��j^a�Q�Z�BU$*"z��[f���@���XC%�KW�f�B��8m~K��s�7����P*$�?;pHF�QV��cۡd�=�`k^ٶ\�>�̀����C������(�z+A6�4�u]�U(F�D�Q���IѠ��i%
2�m��ϙZ1M��}��]g8TŚ.����߁���f Tm�Ic�^��D$J���7��UŒZ`5D�A��C"��iZ�Җ��S��­������f_r ƴ����Z��Ĉ.�5�(1��"��
P���׫���t]'��1�k�1�_�D��2�YC�h*���a}�r=r�&�b(eYs�<6��n�D �Rҙ]��S�O�:�2 �;9���>YP]P���)�&nE��Rh�"�Eg�ΑBY� �d"��fn&���;$322�2�ڮ���ؾ��O~��?��ĸX���`��Y�������.Ʀk�1�[t- X���Ņ[_����f��'�����]�Q���޽{�֭�����˯������sbft��$,�uI?5{	5J��Ab�|U�uׅ�B���ّ�Q]�3B�l�Z#̀= b�`Tu��!$D��ع8�)�|���u�|����(����8����J�V\�ʶ����%����^��Y�	��y͓���y 5��vQ�R%RT�B@�;t�*I�'j��u�!�9�pb���mq�Td�����*t]!����z@,N��gA�� h� �.�� ECr�(�L�	�e�BUc�v��b�D)�Q�k#0Qr#VU F"���C)5�����9%&2)��Q`Z ��9��!�i�
F�@��)5�h>oT%����!a:��C *DT��;/��4{�'���_b�Ƃ!*�Q�r�b�H��*B��{"6�%D  Q(� �Ϝh���(�X�̒31���	�!�j��b��Q��a���V�������A�d�Z��cWyo�������VF"�Ԋ�i������-D<;?�8�0���М-Z�f��>�F¿��ue>�Rs������T#�~��5�R�|/�rj OFu]/��bᘈ �D��i@�h��I�����*�����=9 �	��� ����+67&E�bd���B{�V{X�����Z���uf�DU���|�W��� �de��m�&�R��f��.(�4�S&�0����R��<��ϯ�����G{ۣ���e��`�h��7^R���J�b%b`cb��"Ҷ��е]�
�*jCdr���+�%�.AĞSD$��J �A���E�Z��J�@���{nK���LdGQdm��������?��Ow67��;��@��}��;��U���9v]'gg��������h4��s�z�s�$89=���&�ڶ	Q��ַ����}������U������(H��-6��e=k�5�c!��M�I"Q��x2�׆��uFu]�u��t�v]��(�c&��Ļ�`��f睫�К
w*N� $%U-;��m5���[SuF����A��6%�NW�j�MZ�&�U5��#a�q6����v�w(;�l�`y��uY���,�`�=��>��q $F4�PŢ�	�"��y[ʷ���UJfgz��g9b����XM<""�����! b�1qQ�p�o��'�O���y�|��k�<�fU�A�2nU!h]����s(�8�1�Qq�ci�3 �(a*�g���1"�ȏ��2d����6�TUB��*h���iD�B������MM�"��v�X�1�8�T��xԐ��|>;��/rTUZ�b�`�^�w�cC B�+��(wbef�1�4�p��r{vN�!Ɛ�u5�wЁ��Lh�0h�&����`�vQiCW\4bB����Q<Ѣ�c�� �8	&��G�լ���8�B7��C�Z:�/���,�.�IT�jww�G?����z�6������O�>E��C"J�t�������k��{_7��.Ӏ��j�р�$�p��љ����]|b�A������8��y����nm����_��W����=u��ǔ����Q	m\:���Mp�z��u�, �D��4�`�m �9��b��EB���9Vާ�m%\��u�I%�VVW����w�ȳgϞ>yֶ��6H�c�嬍�,�����Y�r�����D[�"��aJ���Kqsp�����R̔¦l� '3��(0�4�(�]��zSr�&���c1D��뺺� '	@	�.~�yq��L���X�M�4�[����?>���v~eee<��ͦ��}]�+��������!��]�_�f�I=�G����۷o߾]U���b}c�9��:�m��;;;�[�k������W�����>>>�!�!\2%C�
W��&��	�m�v�m�ީ�?>:z���&�b�d��d��b,u��說bf�ˢe��RGP��*!r�($F��n>�[�=���Ё'��B@��%t�a	�]dе�� 1/=7�k�h����Uu}���m����3��b���^	Y$?5�AN��r�G�m��y�hcF�$�e���)F����
��*��$&��%Q�r��n��[�<Fxdj��w+0MBt������ޞ�Ƴ������眛喵GH�A$������U�ʇ���Y ?o�Ւ�lPDt������:�z��`,=!O% �2#�V����"R;N��Ľ՗e]���bd����90"W�-dl.Uj[Y�Z�Z�C4z;b��g !flUb�ʝ8 ��w��'�����x )
 ��t޶��Ԯ��|����3 `b�<�����97OF��#.�,��l�K����~���>�&α���L���~�feVL�@���
 (r�6'�|Ś1�䇥u ��i�sԻ�,��k�M�Q]�U�4Dr̖_*Q�+�%���Ţi[��L����	��WM�)bĸ������t������Ӌ��{��?<===:>�|UJqa ��c(凫��V�,��|��R�*e��c4��$Ƕds����U	�Qؿ��i�9��������xpt�{����?��?��?�|���4����#��F3�P(����_K���k���Q�K�!'�'�0t��.,��뺮kͲ4W ���u��-���|$���Qd4}��G��������_}�QK��u���(���M����5�L��>p��%�m�<ךy1�9��.�����$��0�%j,2��|(!	�(�zi�
�1�y�u �f4�YBH)��i���]l���[�����xur��;�g�'��O�y�j��Ǐ�NO���ַ�n����?]����Y��?x��%(L�����x<:9=���G����[׮�Ǉ�''�;[򣍝:��4�9�+�hx�%��6��4m�"���'?�)0V�#���/�~�u��Gf�Ii��`���B�d�F4�@������|6�Bl��%GU9�fW�1Z�)^y�ޫA��"b4	%*h"@�D�d�1W������f�4ι��?�я��qӴ�o���o>��eD�#�2�=������0?���kn�QU��� j?�/��~^�-S�	
NQ��̚5���Mh4�BXs^���iM��L,*!�#3߹����ú���vw��_|�E�4�;�E��n�5�T�P<^�{�&~��2��jmA��(Q-��um�61!h�5?�����'��H����$ќ��	���}J�BE5�`Dtc�r����A �\�x���B�}gTA$ZW8�G͘NͧC�����٦�ǄU�V��VWV'�����v�s�5m�`����u;f�F H�#�Γ�̮v���""�c���T�F�Db��Ȅ�
�׬�!���b] �:~iI��$����wh(�P�?�ɜD
D�����D��*W�B*-*Z6��[*�uexRQDC�#qi����c�[[[�w�|��g������|6�N���������g����ZEK&spv��}�p���<P@��d��O*��1=q탩*؎��``��ewm8em�nnm����m��������~��_�/�����?����W]�1�X�q��� �F��>I���ߖ����+� `��hD�!����%�?�(!J��]Rr4��TV��v+)�� ��"w��y��wON���W�Զ������=|xz|�����˯;(R�MBn�1�ԧ2�m	J^a�-R@�h�Ւo� �
�2
LJ�<����a`RL�m�u'�����[[�\AP���Ft]0�	 �=*$k[�i���ʶ+3Ҁ��$��9�+Ｙd�53��_}$[�����������r�嫗_���W�^�>8<9?���;��?x��իW������Ţ=o.�?.Qvwn���ӝ[۷��>��ժ��Q@�y��7���;��n�u���_��l6��꒘��	�ϗN.�FE�j����?��O���o���b����/���|���9y��9�뺪<3a]��y>츳2SJ!�B�vU��wmq<��9�
��e��j4I�@&K��Y� dc���*'�o����D|��'��`oo﷿�b{{������Ï$���Q���=�mXF���o�ߥ)��u�� ZT�l� �E�# J�),��XWe�(�5C�\�EZ1
���=�uhC��vۻ�}�a׵�w�
?��wvw�NO_�x.�ک�%;Y�c�
Pc�T�W�yV��)���D�h}������*"l�f6�v��+���m��O�7�O�zKO��+�*���H� D�����0PLuLB*������P�O�"D�΁B��Q�1iI�ڇ��
��Hh�E�-l{�����DTAq4�0�d\;_ҢY4��C(�g ��X�  ���rx_�U]�+��cWb`�ZR#���S�0��
�E3Z�ℑ�œk���F$�H��  �j3�dB�����9v�u��P�3сU�@��}a�����A4Ġ1�UUW5 t]bT�.f6�����'�b�v������
�Y���*{U����B:�B@Ī���e����en����|9DSx��b|_���/#���,{�7�K������ �Dl�v<o��<~���'O.����^;v��h>���
!(!{s�MH:~�9,�c��e��g�����R�˪3r�D	" 2������)B���Ѯpaf@@�)�\ՒE��d��erm�.�������/~����g����?��/�w����~���%?D�1�n�z���>��ͦ셝�G>h�d���@���Sڴ����!�@�g���Ǿ�s�����4���\���b숼B�!���b���b���#!Z:{NI�Y019�(#��;� D�Q�J��Z�u>���v*�����+++Q����/>����㓓��Sh�N	^�z������,�<��4�Np}ss�h��x�s���;���\��Q��_}����W{�������������m��xD��,���n\=� �L�6�뫫k���_��_�U�QE��������_�*1YFi���v!v]�
jI#�{�}�ӥ���%�ѱ�Ω��DY%�:�,?W�s������5scJ""�����`���C/1{>'��{���ʃD���������ޝ{ι���޽sv~օHޙ�MX.O����Fn�(��������>��djg{px� 1Q*����R���*-��b���TAUԥ�0lmmooo��?���O�]UU���ޏwn��{����,��|�F)E�D"���B�-E�D��BS �%�Y�	��FQ�~���Tq_�A��c���ڗ2�"Q5F��#��Yf��S&���Z7KDdE� �4�%�R�MՔ�K�KUU��Qر�u�.Dk�KH�ι�ֶmc1�H�}� ������@�E��d�=�� �S1HE�rA}�HdZ��������<3$B�0�>�(:f�"�A@m?_5�3�#tK��������B��moX�ESרL�ެL��*-6��(
� zq~�����h��ի�Ã���E� b�!�XO���� m�����~c���{�D���iLS�*n ���������'����*z~v�"ȄH1�W�pYC�b��s�, �.fe��
+�*jxT�t<���g��_�w�sv�QTQI�y��tE���|:�޹{��>�����O~���������BD$�2�������/Ib�/�/���xr��H/_�F/w�N��i����<�0��@ �>�J���TR�u���1!�F���d%�3;1XR|�E��? tm��[wv���ܹ�7��;�7v�.�!��%�����_��ϯNn_�T�k�_m��׃":"B�6�斈0�ܔ�����/E]Ɍ��6���Úg� ]��uI���~BM]�A2]hv[��H
���� �=Ē��p��3t	�ȯu�}`$�6��b��㯿������+�k�G�m���ٗ_~�����'g'���qxx%���=��	a��2^�|�ч���M�[����Zߜ|���_�����>����ޟ���/��;��ww�Y׵�t-=g�/��7&m����x���5���Y�R�5�h4�H5;k��lX�sl�b�
-  �Z%�miB4����sU]ŮcF"@"
�z��JC�"��{k\s]֥Y����1FY,�kk�[[[��o�Gc"�n1�7m%9,���2L�d�)J.?F?5�`�S�5f&���6,<|y�(g�Y�*�q�2b
UĄ�%+�%����h/v�`������l�VUoݺ�ރGmیFc�}�Xq"�ɶ�ŀ���c7��fBwv֞��¨���D+�*q�T�+]۶m��nn?`��k�IL5�����Y��s���CTB�h](C���i BTQU	j�{ʂXBO}�� �R!�@$D4M��%ABr�U"1$Z��!h�u��P��HE		��3��.�J�	 ��șV�L诹qV�q�v6:�L�ѱ�Ԓ�h~���C����8j������@�R�t)���/^� H��?	82�]H��� ���K^uB��RUUgg'�W�E�kۨ�������u]�u���,�*U=�L&�|qpx�4�����t����9RX�a����W��d4>9>��7����������ƣ�/�����b��Ѣ=��+�[@~��aG05��(�76o6'��l6۠�~|�)�Z��[�@�Z ޻����������'��?����������/����:��".a��~G��RC�+�bz��B�����;���=�OC�^���TK��5[D@,���C��f_|�����x<^]]}����OOOC�=V��ȑs.����w���G�M&�ܽ;w_�z�����W^���<56V�e4�F�&��cf��B�����:����/8߮����������o��1��aQ1Jn�yݴ懑�+�3u�PcX�C�򏉘TT�P��&�A�՘�K�H�h 13�&z���
z3�P��Jb\4v<YY��{��ӹsn:�~��wv��ɟ���ã����/_������&1�{��êv!�����l������_��<z��]�̛E�.>���۷v��W�z��#��������{-� �@2���Ԓj�� ��ӓ����O>�8�ptt�����BВV��!� ��������x4><<<<:����m�Sbj���H��� ����g�}��������ڴ�^g~]����_˫}�Iٔ,38Ϯm��/^޹s�������v=moo���ۋ�����>�IT�wI���$��n�8)?2���L�\�f�2PEʹDQ&�<���~+��r��
Jp�P�� �P��~���޻�"�������x�D�9c4/3���Φ/_�d�ׯ��fc��"2�j3I�H!b��
]8>>�UAb��V%*A�Ryy+����z��lI> j�r1FF&@�e��FI�؈���ڻ
�.ݧ@������+ �xfbk[��%DQb����uB�F���$���^��A��*Qc���w�B k�i���Dd�V��G%$�*&E��Aa�M�)�H�%GD�4�_�0�d7� �,u���U�o	�W�!�cR2=�x���" �N��P"�Q�3��7���dr��m$Z����cgM�E;"�]x������\U жMh[�)%�sxw��V����g�}�4�۷�,��ggG���Dlɽ��E@�]�W�HMȨ�b*�*q�D����i$ @9��4��V��\����c�(�9��k]J4l[���mi
��sl{REƣ�|�|��_������/_���_�x��9gݴa)�������X͘,��>X�j\LH�ʤ/]-��|cfR�����/^$<Rd<�ܽwo{{[UC�Z8���"�1�|�r��^۶S�=�R{�=Q�Ғ�7�^=8<���O�G����K�{��~�����<�9��h8��R��z�c�.da�Cn4�'c�EK�/xvV��e�j2�/16M ��s�.�Lot	1�"@����0[�� ��_OR���R\���U�2q�p����U4t�4+ 8�1Pe"5+�_���)�F}��&�R�Z�I$VUB<??�BC����~����>��O~�?����/^(QM&�W�VWV�l�̻���o������Wn}}������;��WW������]"�����ön9Ť,����}� JF�e\�g�g����'�'?����y���O���+U���D�.t�DE����������ݟ���m���y����x<_��9QD�v"3ף:988|��	!���z��E���; ��u�VV�P���4d_�����s�rͼX�1+�������?��~���^�z�����3��O��(����́�I�i����02ӂ)?�|���C���C` ��TSrj��Lɗ=��ĒD�`Q䕭0 �2
�'"�QC�Ѩ��O?�������-b~���O�>m��9_J�����������{�h�Ngg�g��;w�lln1Q5�ɟ4!\L/��Y7�88:z��!�c��ZB��	��WV�J	&B�И8s���c�!
X�
�e�l�����⑜�ĮW���aO$���H	
@)В%	Ҥ���jH�cs(W_���PU%F7��J>Ƙ�n ��S�(��Z��=��J�
���k��CF��%�S�Pi�q�H�@Y��0�è�X5QUUDL@ι��ճ�3c��m�J��Xǽ�K��U�X��Z8H�N��'�����H���$p�
%����#�d���Hd'՚�VU�4�������!t�y��jh,��N
;�Yy�-�$�,�����������a0V��~u^'1�Ң�L̥��R�����_���&�C�����_����_����UU��X���6��P%�_���V�D1=p.� ED� X��1P^�dDK�%bvl�̼��R�F"QE�4��B۴�9kg<�N��K]XR���h,Z��	�(*{�^-����- 89>�8;7;;�x��.�Y���M1��KFy!�Q%�/�%���T���%_Âq鐜;�,c��f�3��㔨���.�O��:�0{�c۶��
��3��2ݒ�D��V��,T��M11��qH)eB@)Ȉ��]�ݎd�"�(y�k�;`�7@�lD��}�z����Dr�qѴ_��|�|��G��������#B���;_�#r<�T��W�<�����?����i����fӋ�Ofm�=|��|��'[���bqvrvzzzqqAuňҧ����I�K��g�{����������i������6M����̋��r�9%��i�9�-�8��U`�,,U���x:�����c���萐�����	679˱4��BD����i��=�,6��U�v�>D�Z)e�" ����/�<::Z[]N�O��/05Y�b!��,�~�V����H�<�4M����%q)^�'-(���-�=9q�F���cp�0ʅs%����  Q|����p���x�֭�x<����ڶ��0�ӂ��2�
�fa�;b��x4��޽wg疕1[����%�i�Y�" "��TB������*�՗_*O�jNT0c���,M�9�u@�4��?��	�$���C!ƨ1�L�tlD̖O���mͽ&"U�N�Ƨ��hE�
��ll�1FKٹq1%l$S#iz��*!;ۘ��R(���"M��eG��)���:d�S����H �JTrn{�frU
��E@�{�H]{ �%E���N����K�
FD�kk�&�es8�=�v�0Ep̳�l6�e��(X7@AA�ȳ}�o��]���X�H�6"⽇l ������u�vG TId�
`ܬeJ4��`t�r�W��rr���xi��X�ѬȔu�޺�(��j;B�UU�VV��m�L�3"���t����_U!��hx�GJ��8���L����ZW5Y]��xtp8�N��B@єQy���W����%�1�à����@JJ�����Ĉpvrz|tb��(��������(���(�Aƭ�±�{�XV��X�E��!-���$���������î�f��������ޞ�ez��"F�UԠ�ad �ؚ��s����K�aM1���<�+�cj�f��*��e�Y�R&��F��
�&B*1�b��$K�c���D��LΧ��ǫ��+�m��i��IlBs�ރ��ӕ�vLHUU�G�Q]�ē�O?������2o��?�����W��Ϸn�^�X?:���ɏ�����ώ��s������:��M=[Q��+dz���Ϟգ�Uaeu5�B��@d�f"_W�� �����m�6�(�hy_.J�P���y�P��<Y!�-�QF�oz-���{���2��.����2kE��w1��/_�sbr�9r�
r��D�X�����=\H��` (8}��LC"B ��1%$3�ɤ0�@��&Q���B*�BR)�/�;�{Q%�
��fM/1`9%��@d��tzqq�*� �c��QU�1V�M8ƕɊ���ŹDQ��͌�l�qa>�A��j��6/j(����� .-����k�aD9==�{����ʓ�O&�	���Rv��Y�w�Ȫ�����ġ&�ޮ(�:�˶����`� L̎�P�"1R�L���gߠ����ȱs�;[O�{Ƚk�,QAd{�f^�@�Z�7:x+���b@H�d�$�IR�%ˎ��>�2@Dk�c;�٭��߿��o�y���-,D�RE�]��%�ɞGD�}��(���#jys�<ň��l�ڡ��14ǥ��vkk�ZEAn�DdfYyk�X���YR�j=#��}�!M}�֦� ti)���6[/O�H.I�+�ih���$���C�mqǬ�M�2���:��!XP�z5�=����˙�Y� (,���S�NW�"�s���R��� ����9�`n~�J���Ĩ/�Hc�:_�l�$en~#�eI�������R��4�����r
*H(�ֆ.]�
Ev�uҶ�����������>��L�����z� KC{�%tbc�
L�c�B�zY��J�b�>-7�������H�\�q�PJv�Q�1"W�mBv���mA"Ոy?p��a���׷��v�J�M���̣�p�X4Ӷݢk�N��_l�����#&�16M#Q�������{�����lss�����o��޽�+���ǟN/vw�����˿���{{U]�#L�/7���B4er�'"	�1�H]��hd �gfj۶�1�V�o	1�y��������S"
1���g�b�*3���n#fI��^���:KHP��7ٔ�I��qH�"���]������w`Y��|m�6d�1}<\p0�'���B`^DR=,@F*
z�lG`T@��R�W4�i�mS��ߘMʴnb��d����C�ޫh:��y�z�%�(3`�����E���cx��g��f23��؀p�*��"Y=v*MS�B���QQ�
�G�\�	PD:=;]4����x,�F0A	 �(��L��cI$��4���i���j�/:xk�ӳ����{���~�ʲ	��#$�j�:"�&?MVUb����Pi6жm�6++�F y�<GL�S ��&_�P�BD��;�@b#�����]���rQEN�H�0��9��V�&?����˗/��b4���Cx8;��}��m�9��"p̆+���-�v���WEK�2S �^[�1�̃v́�]���
����Y�%I���������Fd,�DfVeeVu-]t!B����!#����<)�/�3(2�`x
�d�.���kϪ�*#2c�q�{���f�:j���]"2��̈{��q77SS���O��[k���k�Sf�?�N�
݋��Z$��%Q,5B����Do�V�q�<��Ei3nWHb��g��1F ��ט�>U�-���1!Jq��I�u��	�������ߏ�E(
U��d�,i��T��a\��4-'"k��bjҚ��.=8w�K�(����`�Eе�Z���P%O�|��#Q�(��ya��w��1��� "�M�b��@>y��oWF,��`���j0�dW��e��>��\7u]��|.��H�Oܶ���j�7U��N�W���cc�^���{��c����p)�Z)`(����{mZ�,�x�g	ٔ	�izv67�7�Ɵ������������F#c������i5��,	������776�>~��翝ͧEᴾ7���~��|h���$i?�d�^y�o;!Q���z^!bQ��y�} c����
�:�SD�7>p ����X.�(��٩�noI�d3s�>��i�z*,}��ǂ֝��W�.��I&l���s����}ϼ ��;H߱4�Z������|zv��@�UX�*��ڭ!d�T�����+r�cDI5�H���{�4	e��2o��В��:�"QU��5�����$�ȱ	11�o_џTX�B0 ��z*�ґQTQk�S倰u��냃��7o�������Y(��{���(�y����6�� ҕ��M�gυHI�����`w�XX1&$�8Y:��s�`��H�	 kH��HT���4H� ��z-�0�EȲuk���iC�1"��B���D�8��$L
@Z�#9���6��w8\1�ʲ���z��;�
w?�wt|DHZ=JDhS��9���RŜ4]r���Y�.�V��E0%)�b�m ��I)�E_7J��\�۶{GTca�9�:	s�<G�������K���ի�8)z�5'�]���@��C6����/N�4R��+�;�RQ�F,�sO�s�p�d��3��;7d×Y�k�0��;�;D-��7�����OZ\�(�܏.b&z5�A#,����G6�4,���W��z� 9&~&@4�_r�0����������y�k���{2�(�vs�vQ��������ϟWum������{1�N�^�({�٬t�M�lݸ�'��O���NOO��k��_~y���_�ctE�g\��23p�( �7 �� ����Y �y!$mW��%iR!M����q�0K1��r�ys�4�1ƈ* �B�������Uaa�
�Ҏ��G����ټz{um����������lvtt\�;w�D���O��^o���}����;�h���~��飓��۷o���L&��t���b����e����j��e����&����J�*M牦��[�:KA��ܽfTȟ x��S��X��j�C&� ,dE2�{���j���AQ�e�_8Z�B@�n���=�����8��Eb�
mhPѺ�mT�W� �h���H��o��K��EZ�y�������M|���s��!�%ù����_~/�:#"a�\I�z��]#��X~-����7!��(X�{O�$]BD0�а4j��Ȉ�h�Tz�I!,R*�F��QDB`U�Ō�E���K7�Z����yp��p0x��oTU���WWu�aF��p�=��;g92
�j8�Ϩ
�"�QP"pR�A�p�[Hj�%� �����_������H�W�\C����5��9*Ԇ�#GCF�&I�� K�9�R��D�]��t�e�X��!k��QF�U���'��(�rmmu8^�v]D���~����ɣ�G�ǈX�ǅ�G�&Ǳ��%�[�m ������8xE6����׭uU]3��`0U̜����|6S�D�!Fp�(���~P1�M����4��' �(ar1F�i�������F��/E.z=�ϥ!Ru�V��[�2����w��$QL I�</?mٛ�vNkS:�M��}���C������/��"�<����ip�'�\u�/����~����������l>S:}Z<fk=;� �!4F���^ξ]ܫ:?���o�,���0�K����{D�
Z�i\XKH��� ˛o�����lw����bp�D�Q�!D����ߺu�_��������&��J��	S�L�U�z�zh���t6�����ht6>��ǃ~�������� ��{�c�!�����c��s�N& XYY�U9T1��E@4���_X2}�;�l���H��s��h������~��������w�~ۘ����ٳ�h�Ν�U-9p��ܼ�s}mu������/��E୷����}�9����j>�� sLD.��|���)=W�������jWU�Q�4�L!U)���WFf�}�,	��)�
���#�O��\��sQ�3(<vuܛ8h��|��6@�;���z>L�BiS|�����H�����vJZu~��4�;j��(j=k��[�~�*!dHbs�d<B $���l��S8w b� M p4�h_n4EQWUMh|��A9��g3�  �ifTOWс�i�cQ:$B�D��8�Zj����0�?Y!R�כ�g_޿��;�~�[����9>=��������^o4�{"c�!�@m�@ā�'R[ˉ$+���ƨ$)a C��MW�Z�6T�h���<Q����4[D4B��C�l�P]o�=
��r�FA���m��)hYk��9��A�+�-d�����^�ɉѩ#D
�E"*����[eY4M]Uu]��7�񸩼s���Rk�έ�@.uBF�$݊�`sTm}H�Q�t�rdKt��-g���ѵ�׶�wD�=Ƙ�?�|>��^�^G��C��B.Z�4Mc���zUU ��Ūm����H��Ʋ�:gڇ
Qc4~�4#�R+��s~_����#���P�1
��e�P�"^��*�3CWi�G�Yh_�>W� �����;��j9_��&U[\vB�@'��\���߾}�Ef�������&�U�����������G��W�\�'@�f���!9�Jf溩A�(
C�0W"��ɺw��K���w��W��[TZk���(�d]*�n�#@t�����������_������{�"!�~���P�s���������_���q��������r2�����71)�(x��]�1���x8����M��G�Z�qj�Ľ��UK�DDT4ZW���"����Vj�p�<7
 a<��Z�K_cG�D�)�~���V�ւ�޿�Z��76�n\����U%��oc�����$$2���ͦ׮_�u��%��X��������r���Xe%f����,�ѥ���R�;��!ɕQ��E�K���<���U���������)́c�������G���k�y�w���f���J�i��M���`&ý���R�%G�g)<wn�.��t���lYK5�~E�ׅy�%�+f|�	^��W�̽�n�^A����Z��d�����p�`�ː_A����"�5�%m��6Z�
S���A���MD!�����ci:������Ã�k;;��vU�?��ӽ�}@6m�[{��4XE���Q$��| �0�ۺ�Š�P����1D��<=9��Ooݺ������QM�̼����ɓ�t��C�Y��n�z��^��Y����4���u{Z�������֞P���ޟ��s�##9�L��N���+">xf.���C#Y���� H2�;�V����W�Y�y�������c�ˢ� ���}�wVVV�޽����(Jc����(
U�֘�#{�κ�ʪ걨x�\T��2$�C@�#8��#-�x$��z���y��۫���{{���3�A�� =���1wpJc����oݺ%"���ι����������u���칈��>��]^cvl$I�b��Y(�QA�7�9�������G�WEђ�<Wb��ڂ��T�5�)����Ic���b��ۖ05��oP�?g�n�9����]e�C��ZW�y	̞�� f�-5�y��<	��.��cN뽔���͛uU�����k�kϟ?>looooo��œ'��S�+��C�@C��]��k�7���fՋ������׭���D	�$�K��|��Ӌ��p2�$ �(N��@<3;gmQ�u�sc�:�>xԢ�z^y������g�~& eQ���M��,XD���_�����������'��g��'�E�*�I9B�nX��W�w�]��k���`��!(
!���K͓{���������QQ��� D�K-L�&  Ed�zu�7ֆ�!���cc�p0!� J�n������,D�G�������o|hB���y}m�F���?y����"R�d�[�� i�-��<@ �h6	KK
�Yӷ-B�O
�[4QTS0%1�����?��������;�s������WVV�ܹ#"?�����H����7�{_�=aaf�v���{�����4MQ�(2�Lp����U/�}_�%~]���uҴ�hKS���w�}.���Z���,m���h�{��$�PMP�o��tV�I�����ń�i�C{>�I���?a\L$"*66���{��mc�����ZQ��p|x<��+k��n��?8<88�uc5�w�(x/"k�[;;���|^�zM�L'��0�����OOO}�,S��X2��� p|r2�LVW�VV1FB�y�����O?�t��SKF��\>����O
��xܨ�a�!$1�(�9D&D�j�" ��x%��r��A�1�����@���%�Jտd	�<�|���g'2���R�o��0e��Q#Oc-r�V.�� cf,)c�������'O��^ ٕ�QUU���("��@R3�@6I��Z���� �E]���\l�� �I��
���l�ƍ�mD��f�{k��At�ʯQ{��Z@�V���o��ׯ_��iU��~���y��;'''/^<�
��H+Z��v͜�*��T��CeT�������"
��`�=抶�dK�RuC����ϒ�1+��k��C�vq�����Wg8 ��ښ����E@�tۮ6n�P�/��[.�>D��:;�����h�(�~��?9=�ͦ�~9�4��WQ�^5M$Q|�[��p�����G(�+������'�'��/��_��-=�B�C��v2���P�)�z�+�jG�@j�E�۲I�D3G�YkB�1�?W+ެ���1��UUi�2c��b:������������_|Y������������;�c�}����������F��5M���$Cd�A4�ӫ�lFO�|�$I���z̬r6�;<����{��mt�V8b^����w����0yf1�ϟ:gQ%�9G@0A�Eط�!Ѽ��u �"L��Z����i��P�AS�1DG6���j:��߳ot�a�N�@�%Kπ������w��]D<���������o�~������P��TQ!�V����r�~��z�[���ܼykss�W������wީ���/�y[}������ �)I��,�r�O���#���5Fg1Gn��R*ݿ81{oɡ�`ƻxA6m��k�Q{AY���!_��^#-��2DŰ5&:�]����!uTS�/���<MDt������5Cv8Z���!��?4�6MÑ��E��RȢ冈�2���������oTU5�LVWW������(����ދ�_���vw��$A�,�# �Qc�9>::8���U7�w�7o�8=:��������(x���4Z
�5�X��[`m�~�⼼A��A���h���W3���e�VU��ڜ�4�X̓���1t!T91u@�j)���]��r����t��o��/��
#k�"�m|c�(��u]�z= 	!x�cd��;u]7M�EL����c`m)�խ�oT�M}��z�*�q&B����Sg�pe��ݻH��6���1 P�^H���Tx䲳""Xו�f4���ݿ��d2Y[[{��7�󊐜+���/���z��`���,��H�jqL���@B�*�����Ʋ�@�,L��*�2B��{/|�|`��a¯��)1�?�;��:-��d�	��Ⰼ��CףB�j�u�
�t:}����7���z>t���ͦ���e�[]Y���1F��c�V��(�1����έ�7�>����߾s���;���o\�����������/������Bu"3�x8�0�.�J:G@����_�5ҝm]��w>����߾s�γg�~��o����}�O�<��W��F��������_������!��䓏?y���޿v��_~�����o�q�ƍ��O���lo���;O�>���]D89>F�����l:�M����Jk-x��#�jcИ�p�PU�8gC��pLk�D����;�ai�!q�5ϣ�:uUQ��3�D�v0�!%��6�JY}[��sS1��  ZR	�c?Ԇ�H(�k_Us� �[I�$F1������y�ά��'Ӫ���{~txH�d�dY�5e�P�1�R#�ˎ���r ��X7��Xk�!1P��Z���h(�$z:���]��p4����Z�8�̊��j^��ڞg}��?������C$h��֭�EQlnn\��ڏ~���QS�Ʀ&ԝ���^�8�yS�����g��� *��[�Q*+�C��%
&j����K�t��$�
��o[r	�gJ]�^#�6�m?��#x/9�צ0�/%F���g�b��c� bl]�������k�]���]��p8�L& �}={eBx��{ttԦ���5�F!���ʵk����铧�����7�y�B0���_~���.�	�&7M4HEY��1�
��/M��>ݽ��3{�^]U��h[Q��,*�M��
�����B�>��H�J�% �l )�=��)��}���5AB�!h]GZ��z���M>eRb3`@ �%��R� (��+�:����ƐdM�����Z�-iJ+e� D13ks4Ƅ���#�AD��A]Q�Z��f,ԈS��<�;[��X $�,����"RU�(��,f��Ç{��d6�{�~]� ����dG�_뜳N[�u֭��7� ��������ֶs��7�\[[��_L�S�%�HZ� h��۵�n��6��' u%L�[H�Ivr�A�5��P�v�Z�ʌr�u���VY@���y��<�B;�;��*�����ą������G���O�)3�m�< �ob�9���ѣ�l��gggEQ��뺎1���'O��CɄ#h�* dĎA�'���lZ��t6�!Xc���~�_��1�D�dtGQmp$�!���	^8B�/H1z!BR)LA��*��f��j���Ӿj��T$"F��!�몴��������W���~��_|��w���������O�k׮���������O?Y[]�����vm}���}��������?�����������������/�_����{�}��������o>��������?���O��p?��Rzda��?R宔��H֘�?�L���������qAD���_4{��zj��*y%��A��Ϣ(�1�Ʉ�˲,�2+��2M�i^,xx�*]�7�ٿ�"����"آ0��!o���ҍc�7����o��Ư~�aY�w���p4>>��E��-)�Dfac1�5��^ɡY�~�A�`�%Դ�sNa�k�N��}�ɧ����������~����9>={��b4Z�whԆ$
��\̬�ˢ(����ӧ���/����}�{��}���6�Y�F+CW����
�1���U�ѥW:կ8t��N�^~B�/Q�L��=C.��m";�K��y'@�S����w�[�^H�	��G�6|Y@S-�H?i]X����~8���R �)&��ч�Z�4���G �4�����b0���1GCV *W�򗿜�g��g!r�V���PF�&�yU������>;=9��׶�5!E1ϼ_��μ$@���21F ��z"2���er�N����X�����R嘪�ˑ��M�}+Yb�fZ]���D |	����!�	�Q_�Ë�H�,I� 3��������m�DF�Һ��e����d��9����޽�Ec ���D��Aj��졲���̜t(B��(BN$������Z���Q�6 `���Ȃ
e���S{c����h���"Dk��Y{��Y���l6��Q�\E�UUW�9"�z=��h  ��B4&yp��[7o�,�r8ll��țo�9�6��VF+����Ht��r��߹yI$Q$Ԧ���Us�P�~�����:�8�$�;��ݩ&r��DPc�{���R#t�hKv2�Q]�Ż���[���z��R��O�G��󳶑��l	�b`8��l�C���({u]?�}���x|vrr D4�L����,��4���T��>3c����O���o~뽝��{�����o~��`�?::��5- H1Yq���Z��&ɴ㢈�!c�>9�/�v�9�f�.VJ1ƨ��>H�W�f��i�6�n�~meuE�rJW�$�͵�k��&�c��,ʕ�J���t�+ʭͭ��5_7�17���s�|>�ޯ���F���YZ��O�vw�A���Yؠ�!�? EQe�,K�{`JJ ��px6���nll�E9���Y�1&�X�U��b���<�,��4���E��u]纓����Jc�_:��qC�,ED���6��G���"Zn�ݓ� �ykk}4�h|�޷�������h��6�\�ѷ�V7֘��t>�=H
+^�ĻI�s��e���nFBK6����U���j����/>���ް���.3�F��|��NUU8kc� �����F���˲�L�w����7����|o2�|��;=;=::�Ng�n�VF��2����� Xc���E|%R��)��x�8e��L�<�Hx�0m��?ag���ϴ�}��d����X2�N7Bђ��v���W���E�҅b�C��c�!x�N���˩��8k]Q @k ���9C��+��lz|t��[o��{G��+�+�����IY��A�����b�� K�G�&4�Zk���uJ�ʞsf:�%}6���+\]���]�s6�k��@jJ:�{�> �!�.�y)�P%D ��������@��0GH�a���̑�,�E�6],����W$�]�ma�]a�1�#��`񒥢O�^�k�l��. m�(�$c����BE�9F������~�������+M��'�T2�Ǣ5]��X}UȒi B����i���[��ƻκ����(C�O?�L��)��GU����z��7E����p�h�2^�x���WU��R��h4��7��������ݧO���_�x�󕕕w�}w<�̦SѮ�|��z�`��Լ�jXѾ	N��)r��z�n�-*�c�C �*�N�/�4�^�UEZ���5������b�@g���*|�ͮ,v��@ m���1�%���y���B��������t6�!�u�Z+�!xL|8V�յ���p8�͘�,K�ΦuU#&��l6=::6ƾq�������%��|�;k��ɴ��#R�Y��D�#��1I��$"
�Dtֲ����19�#��t�'����?��2/�*�ñ�k�!�>����W�7�������w?���~<�����~:������?���=�?�����������{ιL&�O>�����������/���/����?~��_�OO�c@ ]��HH���|�7�Sͫg�w'���kMjl�������pebh���9|2F��d~�Q=�it��ǩUi��brc"��f/m �,%����m����Hu�Պ@e\Az�����j�s�c<;;���z�k'�'�`�߳�f���'@&5�S?� R�/YS)�O=\�\�ˍsˮy�!*$�\׵+�r�{��Z�^����B"��w I�Y�������Ç�:�e�WD����\����������^��F���w����x�/���ٹ6���o>�����(\]7eQ �:��@�!BS7i�-��bשjWJrS;��o�8�r�y�!5��K�Sfw2��3�]��bl��A��D����i�W�"5㼯��..�K��Pz1� "�{c�6+�hDX�� ŧ$�hmҐ��Դ�"D 96�#��0D�� �l6�M���C8<:<==�ٹ���V�ՃG����9��{��1�@��N"�}����y�,Ε��
BCd�LK�@D0�𥔄��NF	���"3�A@����.OQ�( "Ʈ���;E� ��Q5�Оk��K/xy�)NdȀ�r��s��e�����C��h
2D�Z$�pu\?�s�E��C�$���L�,F&MR����ڐ�-�i���Wf%W!g�!�����;o�F��++ rr2�'�X7M���څ3�J��1[�H��{���۷o����ы��u��o�����D��"�o�.���������λ�������k2,�A_������> fu�C�D��"�̂�©<g�����#���~��_�-��Y�T$Y�o��ӹ��<�guԋ�u��̖����  )�✽���o�mu#z����=��o 2p+����'�4d��u�,׮]{�ͷ��	3onn���G=|T׵���ܺu����*�Ґ���������o��boo6����[y��n���	�b�dA��q� @�=8�K�.=V�����e_!gGX�
�� >a!cV�ó��_�����s48�濽����O�s�����>}�ྰ���w�F`2������Z>�xtt\���9"M��������1���0��s��~������ۯonoWUupx@4Îdt��1�i���V�
76M�	��������r�������N����֐,G���>r�s�'k���LfIj�)����[�"�h���z�0F��8	9��?����8(������Q�A�! iUjJ�SX	H�h�<s�н���║ƹ�sҼ[Srա-�$Joݾu��mc���7�7�y���g�>����٘��ֆ&HY���c-�������o�u'�0�_�q��/����O����dZŭ�7�O&ƚ�ã���F#f����~<��gƐ�97E��몚 �s�b��$�U��=Y;��'�T���D���ݒ D�h}�s�#c��R;� �t�N�<3�����S?�K1�������:�6�UW�B���;w޾�+�������onM��{{{UU#����	��c�]�>V�V�����OOOC�(b���ڍ����p8l��,{އ�͛ ��jmuuss���(���,
IZkCH�1D��*�	`�T������;;��d��e���z9�d�Abn=�P�BQ�6���E�"��F�0G�l�r� !���v����d�@Eam��J�d�Kc��P1����a�8kU=��g����^}��A�T#4��r�������E�� ���@��8R���H��䴼��O�g'u�v�K���cL�~:�Z�8Ffi��{/�bu���!M�A�BU��ں�b��x6[�ͦ!xc�o^]]�����(����������tE�}mg��r�M��1��x���Q���x\7�p0��"a���w8�_�c�jSb1[[m�F�U#�M�XE��bo��-V�ڥ{+EQ��U���｟���z�<'�}��7'�{jD?��@�#���)�XK�"���1�4�}����/C*g�.��;�u9t^��}� ۠��
�����J�f��߶aյc":Ԫ4! ��L��QƜ�,���Ge�2�4�T��pC[mY���9c�S@ψ��'��5R��.+p����!1��YJ?]m�wA����������HHHb�꛻�q�<���[/���G�6�%��� 1�1�Kv�{�S�6�g~t��)^`��$�"���3�3wb�.(�_�5��E�vo)L7�nC������_�-Ě��E_L�_���0Z�?���ΏOo��64�)؟#�&�S��,����].���ҲV~��*<����A�<
Xa?nw:� ��!�I��]�G@Cw�y�&ei]�E���7�V�E���|��o��*ఋt��D|D����w�G�8R���~r��_�i����)b4�G������p"A%�������t^1dX(u�q�<o�i�}D��r��nG��u���d��L�ۅE���+��ӷ����%%�<������IL���wYvH8	��HP�B���\��5�ϯn�z>]|�z�F�p9~��tW��.����^�|c���3yxx�_�z=�ڍ��r`�^�Y����"��G�]�I��Q%�g��z �g�jx���a�9��/1�N�3��\����,a��c�4��y4diT�;;e#B��,�MjyIL({C�6���J��x��D��T�ǜV����lу�܆:ߜ�����
`(QB5��O��mgkk�<m���9���zZ��8� EO嵮\�1�����Ou���><��d������꧶VB��Kͳ�� e�y�' M3E�4[(�����۲�wd��yn��צ�߂,�Z��I)�,���$..Z�NW��*�˵���:���^
4a��p�q1,KOq�ȸkU:��?��b��X�Ե*�ӻ�9�����~���F�����+��ފ���~�j�8P1��xY�n���b��Ƿ�Ubw���u�w�hjlf��
~Ő���ފ:q�*~���8�?�H?�ҍ� X��e1�����3�ʉO]\]���w��9��"�����А�t���+�z�%vs����i�|�����Oz ����
턖|��\�
�T�w�t��ݓ����ƭB���n�ѨoW�{��U��7�ܒ�X�^�K��&�+yZ��]��v�k�n>�B;߄�kQ#�ꝋi���w?���$���^L��_����c�xR?�4��(�9'A#/0G�+�me�T�z������娨��{˷����4����@��!��Q�L�d~A����S�77�z�IX�kO������k�)WWW�C&�;��2Ғ�W����Y,8�"a���LYw)�lN	R!��Y������ ���=8��������C*Kc2�������?Ē3�=o}B��_b��@�0��,�?��v5�ڜ�2Y�s���;�,/?7��V�mm��g�,b�G9u�#XV�c^����Gʫ��T�k��!ճ�k���Eq �-�t{:���T	NA�J�cv{��l���.*��`�����@�m\[`������ʀ�U��qG�����v,�g�:\&B`O�_�-��>���NԄ�����tXSm�J��Ӊ�D-�ƅ��8���*��4�WR	)[�|rC*�1MJq���9�ZqI�8A�(��#g7�"~��8�ü�p"�-|%�4�?������EFI���=�G�a:��g��I%/7w�<���iT���Q;YZ/ ��6�����!˃�qw�4�c�.����UXvk]<�������a�V��0�F����9��ޤY�[~Y[�G�En�7�ݕ��rbݕ��7Or�� �Ј�c^	�_��l�Ń����YZ��%)��z��޻�Տ���(L.80+_�Ww���r�e�������ZKkk:�z���CH�m�k{�>���B��G�n�����>>��K���=r"�꓈�$�����g�p���:ɮ�����t/��:|��"?׺(�� �:K�!�� ɗOhꔏ�U�2�3Հ��r���t/�b:�Qst�����F}��cp�MH���B�vۚ�7�X��{�eW$4����!�:#[���H��}�
3���9"ƽx�^b��$�=���
i�j*��͗	�lo��_��i�=a7�0Bt���𸇂�����`�ccc1�Q�*=I��cf�l�q�u��� ����!�L"�}N~E����2\� ��KM�QvL��dV��S�=�`	�G�G�G��J�O��%����[���؞�&�r媯d%�_z\�In#{��XWic19�hϤ�I3��ٕ�h��RLz�܀��%y���5��|�>o��Jɱ�M�K�'M����ݘ�W��/O��`�8�uu�:?6��%������N5ˋ���.X��P&"|����sG�B��p���Ϫ=��d��ߊ����@��Wˁ��qc5���;��ᲢY��Bۘ��D��ӉWn�v���?w����Y=P����ջ���"P�R��[�O-WҨ2S0.�B����i��Wl{e�����:�?�?��������
�� ��#��9O�E>|U�^�S�}|��_�y�ғ�gT�ac��3ur�������)���E���s��3;�1���-�?s৚�]L��Ћ �A���r;Q��qb�?�ӑ��,c���G�o
�\��sR��l��(t������r�G�
���ˀ-.����[�~���'����<�Ys~��f���\~��4����p$$����LU�s��r|9T�v%�fq�o�6��ѿ��(M=��������	��hhm� �wL��$������v������x�D_]i'$&�����/��{��w��������P��D~� \c�>�Y!E��+�|_�d�k��*�z����@�B�98bsB��[F�]}F͓j�w�O��.����P��W˃o��-/���a[����9\M��O\)�[��^ư)ʃ_Dra2�zDq�E1t
I�'x�C�tt��2TT挘p>D�1�]p�k�����.�Y")=w�]]wd}ӽE�W!��O��D{��s���ߺ�������I�"�I�Be�Y�����dۉ��4!=��=j����^�@�q\b޼�LzD6��5(���A����߄��YJA�Lx��f}�?�_L�7'��'%�*c�̱�m�09H��>���/���0�V������ͥ9�e�u%p�����/������i�E)�Rߟ�LW3@�-�4(M�?~,io�'����ώh�����.ba��¨"DڌѱOw�sŦ��O��<L�qJ_v���"9G2�B�f`s�[K�y�k!v��gx������ٹ����e�D�I������A�C���ղ/�rt ��x�]e��b�[!3i���d)r��a!f�_$d ���'u�p����:'K�̦~�K�~\��#|LU%UR3h� yWc����T[\���ٳ@�b��9Il`�5�� �W���L�ݘ�PǠԉ����^8-�������{"]�3�ٞq������(�W2���:�O�syh��ݽ��K)�����s��<���x��B�ª������~2���f���J��%�ň������\M�ձm誃�1Ē�������E6�nv1GFx�&��lhХ���[��-��bf(s��>�Ӹ����hF�#�,����I�#�6��{VW��00<d�r�����s�:�8F��Ir@�t2I�T׊�CSM�m���F�$+�m��Y�0�	�}�ʫ85�j�Gq����Q�G_c#�׽�h\���(�T���`�Q�g��'��_J.�׏�|�Ē#Ii��^�>�,�",2���:�f2�oe�e
�!a�Env�l������ d�Xp'F!(}yt-7�L���I���i�]/A�۲ߟ����� ���ƫ8��!�`?/�����|��T�2&�b58�ֶ���iA���7R�W�k�����U&��Z�%�?����s&�*D��7�[n�w�'�!��,�;��t��,;ȃY���������{�Η0����F1�3�2�<�}]b/��kv������g G�-#}�r^�ͧ3wtN�o8z��b)h]��8��ڢDK>*�ݶm?k���4<-�M@:l!����!�w
��E�M�bI�#�z���b�'6��EP/�j���C<�͗A����]\\"�w����{�����t����G��.�jl��I�*��JЍɃ��|).ΐ81ܰ��3V�\��ϗy����6kaa�G(�y��`V�����]�wr�p�|"@7C1���R����"�e�P	����w�K�tM2�K�39�.��IF��JWO�����Sn`���yZ����c�j�-}�Ϊ0*����4Y�8����ڌ���.4�c�1:�ػ�o�Fj�:���p�md��<�(N+�l)�7�B�븚�R�:���w���P�� ��rg�kK6�:n.��`�m���4������t�*(X��/A���y����9�/ݚ��\3yta� ](���}���Y���d������넢$g��PE���n>)��A�c;�h�x���['A�ˌ�e����B@V��R|���o� WU����o����&E3c�6��C����`	?'m��qپ��R�̍%}*�}i���/uf����X�2�@x�W�]n��Mt� pgDn�CB��@ �ӿ��t����g-�O�h{4Q��1b�ь��A�칝�_�h2�?�ξ|%���TC��y����y��es�&L�P3�?`[ev��i|�Lb~��ű��mݑ�#*��}�2����.s�̜�7��슊�]h����<�[�����n韛3�Ҟ��F��?�M��*�u+�!S��s��.�� :���D��=<7;��+Q�/����"EN%	�OJ���"�J������ �K�W��Ĵ(�L��~���sЈ�P�U<}��W���rU�~o��*�BWw�6?,�����E�P�b_80�|����E'�I	Z%��l�ğ�Slj�*�L���k���H=�t���g:�����C;����(6���fbr�3���曰�Jۃx	����`�/�U-�m�[�[h\��o류;켛�>?M]g}B7jl4�+�}��ƈ��x��T�i֞
���u���1����]����Ж%ea�!/�"FoCh���G��׫B@�0LE�r��p�'����xϸ�b�����}I���/Y=��5/6���M���>�
A)�ӊ	c�A])���Ua$n-�!�k��A`�ƅە.~�ƫ�s�б�v	)z��_�$�ƶ��yG��a,������r����?����+~���G�[�3�3���t5i�'��þ����110>}��s��i0��}h<�CV�`!�Ѕ�h�.Ǵ�	��ъ���F���97;�ER*%5Rt�~�IPiΊ( ��z��ˤaz[a�M YD�;l!`�W[��@�uzEӷ���;�U��e��eMQ[^ ��7�3,��2�&6�T����T�b.;�F�+��8≇��G<���t~RR
Aa�|�����6�p�`F��u5L�j΀�{�E?R�$ (R�~���9C��o�2KK��]]ߎHQ���'cn�7++�ssP�[��������sQ�l(@��z8�E��K��u��L4�=� ��翎u(��SB��%-���La���<b��3�
�� 1\�m>
L=�7�ݰ�ʎ�# �\��#16\ϡD�S1�$�lh���\U�7�yHQ ���$wa�fi��`��05�g����o��B�hXv����?3)~ ��(ңD%�%)�z�e���|;�<�6��S[�o@@����q)���߭��Ƽ`
E�vn�� ,;[߇��,,gD64ߛ�����c�4j9��.���q��Sě�Qv~�M��X��x@��(�sN���D��8��?�RY;>�QYr�:�� ����C�ſ]�
��Fs��w�Ǎ���*j�QsPꇉ��P�B���EO�,.���Ë����N�D�BH��3#�X��cn���z���t�C�K�dYszX��X�`�ϟ��O�5◍�:�
�e�$k��$���ޗ�ln(�+�|$�&!�4l��p
Ҫ	�>����3��d���XoڣWr�Dd��vW�3^m��;0
~i���u*�X��|������!���1{�{��{����>��A��#��7�v{.��}1i5�XI0���F<��y�Z�\(�����s�zEG�4\<���>����%KE���~\s4��⥂�R��-�>����H2k��\�Vv	���%�(��s�/���u��M����>�M��|���LĂ�6�.�S܂�Mx#��}b-�j!���F.w\<P���^F�����.1D沈k��~|����e��ٮ�q�8��g�<w��0�J;r���ͭ�6;=�	�+$�5�P���3�]��oi�iQMC�R�C�¥MJކ��=��\�D8E+�����s�1B�k����蔬������<�uDVXISK�e�8����ϱKb[%*�4{�Fu�Fވ�ts��㚞�W�F��#����0=*<eQ�d�w`#��V�`|��AHh�+- p�#�JB;�t�e<�=ZX���(pYؘ?�D��<�46KImH�9�Q>VҜ|��^�-ilB�[�,|Du}���b	O,�q�C6��B�1{�7��W3b޿k�Y��<����߽2r�����G��Ąoo��Eq���Ԥ�Z~x,�/U����'{����GTO���T�o��p/�����$�����͐���ɩ�(kx����;�j�IN)�"��R���K��?��,����fh�훒�Z<�s�&[>�Nu�³ibTކ���,�pXHr��ZY�h�8� ��� EB������屳���}���Ae�9��u�P��Cշ]�Y�Tg\*������E�zZ}zg��<����%x�O�U@���LAA~.۸[�<w3��<>0y=�U�y]y	&;��=<L�s�9���S)ƉĻـW�@�P�AH�a�C���Y�ՓZ7�	��쿗�" ���]/Is�f��>LP�wʊ�&T�F������g��S��a�Y�,rI��)#��i(,�����<�I��S��;�6Z��X3<c�(N����`<2cP6�~B%��`]�G�gc֮�dz�Z����Z8�vR,q�5�T{����s��3j�:��
W_I��)�<|Ҽ�2�ۍ����w���������_�]^^��\CuҪ�L���r�_��-�+'�K
giT�B*��W�"�PI�BE�v�sk�L��c�w�]�L:;:�Dr��|��Z����gm��$�vζ��yO(*�����=I�K���zV�:�}��B(|�!��#-�+��^�>������.e"!�ځ�d�����,a�t���9�v/D5�s���7&��0���	-m�ԡ�����އV9?7�r�K�8|I^��h$�+��
�z���lc`�]?�އ�u|�Y! �I�*`@���[\�8�l�{����z@U�BC����T�����*>���	���?��J�(Ի�Ub�c�����~�y�Kn���BQH����"X���6_�6)q��Cꉭ���h@�n�wS!A���^�oGd�9�M���$������V'�g�9R2g�t�!��Wϣn�q�JG��BsF�����Ftxm"Z�Gm��"��S��wSˇ�k��<D�Zn~�ި�}t�`o�~r8co�c��I���6��+��\Ϲ���V�of�U���U����j<q[rP�����֊��&�}d߫V'�]�=�1ϴ8�JQ����]$����0U�W�2c�`�L���Z�ea�{­P� YхL�K0A@�;�&k@�h�tCRf8
�{A��߻�Д���ǈh��b���
&-�ݎ�h4-��2��o�y�/�3�(��0�֑�/�P��t_���1�h�L��fR��"� l�B�!V�֧_��4�0x���^@qa^��b��y;�P��5B* ���0ܦ9�~�ϭF<KC��2u{�� /Os�	x|�S�a�9��p|D�7`��nwwU�I���X'�D΄�����[�UV}���7*�G�n�)_�K�Ҏj\��^�L�ff	|�,���)E	�	� ��?�U9��\���z,l�42���޼�aÞ��l�����8㑢�*E㹠|�vW��fy���v��0x���I;I��J��06`�]+� �bi��C�<�>䋟�'%�`&.� SA��р��ۣ� ??����ߏz�n�}E�#��F�������
5q�Ob�ߠ�������ad ��F�^2�	�6��_�.t0�<�:-��ܹg�#�����y��6�WkQ֌����;3>y��PtC�*����F�6
1VY� �����Qv=�`�D����B����V�jaf"2�A�B�O��Qq�>��4b�x][���Y�@dg�B�5ӻ@&���l��@��C��͞�L1�
m�2H(���𼦏E�q��R4ʂ �T�	��т�5U�I}�Ԟʯ)>�Zƽ�ц��+�U�TV!\`ѕy�hW��Q������뒤V���|K�a���g�&��� ��0`l�ɂ��<�Ʊު�6:�w��q<(�����~������R�$5�Ռxܳ�'�D�Y�^��}^}�{�Ǎ1^TS�����'�jg�d��E�%/KҴ ��~Ă�o؋���9� �� �jm-L�穵��^�i*+q��l��[��	P���޿ h9=<'!{݈\Xt�,̀	����n�F��~|Xr&tS�$�mU��uA}l-�-��;r��)d�[[�ܣ772�x�Il������;_J��
٘ꄓE�GV�~m��}\���H�L��"z�f�e%�� �&Q��첖�yYb]DŇ'*:�����ZSW1F�����1;q8�674ۗ'��B�F�$����K�|�?+�Y�@��_��� C���]j$���fɴ�� �a���X�i9��8J�#e]E��$�LI"���+貒��5D�l��<��L�����
�҇��s��<�)l{�8�b�a%��u�7c�$�y]�B塺��T�稟/�,�w��]?`���cӫ����bQI�g�ZK9F�9*j}�����M��������d�m~�F�<����{Vc+�$��Q�H[s�W�Q˩�C�E,I�
��e�e|&�Gb�q���):�ۺ��������#W}����k��n&��=]j��&��ӓI�f���_�R���R��8��pk�X]՘�t�o��Pk0%��TfB���+���xuwKz�����B��	����Pe=�+-]��}2 ����t�mY�:����>��&Qԡ�ޱ�9~�w�c�y�(�E�HE�&%̵��Ɲ,�`В
?�h^�P��{h{p����RѬ�{��wkq��	ɣ0�J.�����hn�!�_�L��1�$�R�3���?.?�v��|�o�-7B�B ,��&�e�$��b�-q��� J`5��P��[p�����Q2���Ox�'xIՊ��pK�y9
,�M$���%���*�SD-7 ݍ1b�;�o�{���w���ϛ��0P����M\�A����{Y`�puɏؗ���k�Y��LU��{�菤��.O���5�sȠ�Z��"˪��e�^��]E�G�:3��M_I���o3^�O�I.K���t9�M��&�6���>-�E�A�(ݟŃa���J��h�|53��\�,��'��� �ǻ��6cAs+D� b�m9b��8��2���L8��|%`w�,��_	�B�"YN>)��܁�1�i7�!n(>�s�n ����z�BE�;m��0v!����6�!K��O�g��Gz���3�nv�O^MI�K{R�5t��f���M��!�X��<3���sey���3{��a@�>a��Ut�4�HoX�<�@f@�pP��fwu�3�yFX�����e�\@Ϫz< 8���{�E����@v��S�\��-��j��5,�)<z�}?$�@T�DP�b�Îr�l��D�����$┈F QN�h�PN�Z'd;7���C3���Z�������_�<�:|�K��s¥��?o^�Ƽ�zW>-0�1�k ebC��ͥv��W��5�&��&`��E#�<E�O&�x�h�Y;$������# f�{JF�p�B_Sa2A�	���y㙬�65o0������'v<q�q��ffP#@���k'z�Of@�O#��O<�ߦ��͚gL��`�T 2����o#fV+��Əs�"����Ӿ�"Z3�OUV�6�wi�lwFUH�dl����BǪg����DW�B��s~��>�W"4@�p�pÕ2�_��,G@8��tx��@�5�۳�G-��:�N�-j�����xy��w�%~�y]Ӹ�ğ�#f�pHɆ`���*X��x�U���Vd�;��Ikyb'�$�K�-B�+44�?�#�8�iO��G͆�W=p6j�}����2�]r������'2���y&�DX�%k��F�u����89u@��6l*oS�g�
(h��-��"( N������� ��	np��E�h���ǰՇh�&�Ю�q%�J�GB�����Iq�l6qk ���I�	B�㣃�_���4�����6��!�O������I�;߳��~�޿����A�뚔�{����{n���k�� /T�k{z���C�+.�j�#�R���s�ϛ��8�,�0BJ����^D�D\6�`cuױ��R�F���>[�8H݆7���;q��ZVhRh(t�����H�H�F
�������݀���a}:�?�8��`��f��s�2*���xa.n�����T9�(���߅	��K�M�ږ�>TLZ�^o��`��H��uѧ��k�G*)�@�މmOj>S2���
�QV�ŵ�������*�7:T�
�i��x�h_�<�Ra���,���fo!	)ii��� �MJT�N6��N�qR-10�SU���1��1�C[��X�,�2�4�7
Gb⼃�Đ���VvI��������_^n0�f�:6�����p&���tL�������"�U�<)�S`�J�R�'T�ҳ+�QSQQ��:�	�"��N���hJ�w���1�ĄE���|/��	P��Xp!
, �N�O�,D����:m�Ca�6�^X�y�RB�/�6���Et���O�S�Ѩ�Ƕ3�� Ն���q[~U��Mˤآ0����Jn�6s��:����N2D��k����<3�qx���s�4/>[Ě�,��و��9���KBe�Y*�I�^n*�q"����X*��}�aBt&Wc�����Um�S'���*��̴���)���%'㕢�	���V5�:1Etu5��]e�b�i����}N��N�X�&!dd�D��\1��uq�B�����B��/m�8�KP�h����e�r��Yw�xYy���@��|ܳ�XlyCҲ���oxve�$	*�����^�o�H�|g�|ݬ�x�,.��1E(K �v��(r|Γ����jwvʉ�Mx�v��R�?{���(�bU�\�ԋ�O@` X��]���3F�w�[��}��=9��π«�N��^t������A�H[.�#��9���ϓ�kM�;��C"q��T�la��8�HT�[�ѽ��U{����o�4��;mʈ�I�`zD�W
�"���e��Q���jC�V2H�����
`8��_вV�$�������a����.M9'��"���HXn���t����H�(:͝�p��-�;԰
�I�Yw�+@:�(Um4��'�\���giO^����>��$nl!5�#��f8YE��	�k#^!N@��c�2���OzT�P��F7Ƕ��6y�*T��ed���V��m�{�G�,W����-����r;y6�w�N��6�p]٥���y�����=�,}�gm���YZ]y��Ȥ��ZtLc��kάRJ���y8D�IH�!%O0|2K�����O��	�q���_v؏�T�;#%1�����1&%{F�rH�c~>�|���˥�
��Ĉn���̫ _�\�&T�. C�`�XmSij��sǛ�'�B�y�E+�����*��1������w�g�d�0e��{��Ao0�eN�&q�>�:�
��� �ڭ�.f� D����E9�~���,3���B�܌��}��/� I<��.]J�By;�z��~\��*��Za��*��"UÁ5���7W^�����*hZ��Ѥ�)t;~�h�g��5n?H�#3�ǦNfl�$i��p�g�y�y��A�t�x\B@�J
�0����_s*	�����}��bQ	発������).)���&Bˍ<Ϩ�zR��Ȧ�A2+��A��I�ﳆ�|��Ϛ{�
G!���KV�)�zr�H�������<U���3p2k�w��&&}E���N�%ڦn˷ed�i�8H����pNS�xO���b&<�������g�nFY�ߩ�Bz����[4�N�j���x���M��{�#�[OPP�������f�}P�=��w��`�W�[pJ3uh���]A+S�h��V%��P���w�)�΁3\H��&P	�����+�h����p����TLj�y���*׳n5h�X�`,p�|}!V[��
ũ��a�ڰ��1�����9��ۆB�mW��[�ed�a�����y�s�qs a!�y�2$Y���2~�f�":�-oݍ�j�����}���"[?YX�6�Y��B����p�8�d��5�o4	LM�A�l^����4']����ۿ�C�d�`�xsv�ǓD}+��^Z��H��^�#-|߶7پ����E�"�+�bJ���f���m��Ŷ�s���y���n�v8�M������D26�@Bԝ����_k����Ж
nA޼~=u����*T�Q[�-���HK!�hM��<;G-k�O�׎jT�q	�es�( �$��]g�{&��]b��6���j��~��^���"��9��~/�5#C�p�x䜦��>Oft�AVE��Tcڇ$�	%8Bv�i�>���g�N�O��y���)0��]%��;*�W��7<�Odx�K���0�"�~mh�?��}�o��+P��,��sL`?[/9ݪ����J�_��
F�*3�#�����e�s��eF~��,G�nhv�7�Vc�VBX�:��V ��11���pi%�ˬ�z�+�Q�rH`ۥ��4P%L�K�z�p9��Q|�[I��hF��������jl�k�
�J�ZaRQ`ׯ���;
����W�����X��� ����Y&7�N�܆�Oՙ���7��bh-���3�SU�l�T_�3�~n�#k�V�-�<�B�A��F�87��������~�~�mh-u�q�)X�!�>@9#L��u8(w+�b��}p5sL4&�f�.�ޖ�gg�Q�=�������9Cd�f��3���TR� u�5Ȧ��Bx�=�#S�#�J���s��QUUUo-nO�g��}a���Ӯ��# ��=V8(������g;qS�F��-,����6����H(�h����K�l;q�⇮���x�)Z�]��(���9���1=e�j�V���v���� Y�S[b����M5�[g^��)�����S����f|�W�����Q�AP@�$NO֞ZHI�O9��Qr�����	�Y������jY��-0�d0�5^�?
����ks�5O�	�[ܯ�4� :��}!l��y=.�1b7@M��~�;���C�����Ҿ�4_l"��uѝQE�VN|Hk�g���N�M'�7Ht3C��Ij}m^�No��E�s��� �f8�E�@5]�f��v��yЗ�7pO6��R
Y�T���>����u謖Y�Mv�.�H&'nl�s�;a_7o9���ٌON�fc�Yّ�z>�ծ)>�n�#�C�\�s��t�N�^Y�����_t,�55.���:@6^�Jc��:��	w�҂�OU����+�6�Ha>A�E1.1y��E�2bR�bkNd�,n�ߑ�wIu��̫�'ψ��v..5��#\#؟���Y |����u�)�zW�XY����Ɔs��7�O~�܅�r�n��c|]��9Ryx͜)N!��H�2k<���&
�������Y���x���F�:֮o�)fm�l"*\P��h����4��o��N��i*ѣ2�L�zgG5�:�k�}�S�x�;s���69/���I�fh	7 �����H Џ@5��u�FlO��Xvlƶ��M�lؾ��͵��hނ���ֈ?��1Q�i_Lږ}M��Ab�fA}�\�7�lH��ʢ�� �� ���To���9�PwO�e���{#�B�!�N�k_�.�m'�p~t�D��]�^ܚ��m��Z�8��3���Ɇ�洺����(w���dt1�_����m,88:�9��z�X9�@:0 �rF*�sy��ʩ=7?�tsp�s{<Ŋ{yxt��<�u3��u]m!�\o���&&&�-�#���8��|�����6�\^�gD�G�H��u��ͤgg�w�q�sM�
=�\�gP�?ŕÿ�-��"2�GP��oG���T����sNy�93:q�B6S��������;��TO��T�M�n"M����_��%#��7i,��G�^젋s?	��k��Q�s>�6�.΀&(�J���@�ǒ BDyZv��a�1E��I�`�&I:�s��O *�y:˿��7r�et�~���G�L]	;X6%��_�<N&�t\~3�~�d%+!v���^��l�q�K*{��a����Mj�a�U1_�t����y�, t����	 F4�OǬ�#Ma�"��
^�u���h;���jѕ,j3>f��k���q��x)��A�u뵝�f&��B)*����q��I���>��x�s��� �F��@rq�-Ta��6�L��CITWC]i(��f���)�v��\��B��^�M*��Q����$��h�8��
�ƕ�g32�5a�x����Ԡ�P��EՖ�r�4P�����s�ܥ��6�P�q��.93���1o�t��21	Ua�$l�P�
mY�n��P��2�>�7�qN��m �?\�Y7��qa�xfQ��Tl��`I�#,�|5jr	� S�h���Z��9��Sr�t=���n
��y�)�gD �W�*#�W������2��0��U�X͚���.��g�{��*-��nxg�R����Mm�l�����G�^�|mr'�)�,�|\�cS𶓸��3�M����'��A�ݮC$�,Eh��p�ˣbXm�ŢV
�fKG����bn��ʕ�՜?�0Ԯ�zt��n�Ӌii���GE�MY
��^-O�u_��[{
�RB�{@�9����m'�yru�r��n�����+gɃ�EX�
t0��Jy�W��r=�����p!�6�D|�JE�I��<H��}�������h�q��8�0�	�����O'��cɫ��ـ�g�(J��xwKoޑe�l&>�[�P����~B�R
���]�R}hy/N�A%4G>{��Cv�Ս�mȳ�kǒ��z�����U~�����K%�u��jC��x���1�;�9B.ޔ��LSR/���P��*�A�Z:��������HmG�7��f
�%�<=�-Ő��d"�A�~�������Wc
��snaH�q�$���"��{��KW��VO�9)ul�Ԋ�W���za�B�X�l��`��Zې�ϝ�������4.��HZ6����Օj��?[+�te�����!Mƥ�2�L�#��7ő�g�Xt�\����1�Zb��ݳ���!��7w��<�B-���&T|�*�0�Nl�{�_��^�$>���#9�w�M)��);�0��j��}�!����_/(��������wr�刺��r��,,tf��x��c�'�lgt�M;��K�O[�g)<���VL�؞��X8$�*����s_cs6��k4��X�=bh���9�	se3��j⊛Nvj-n�2P*f� �/�'�O-Q Ȁ4�u���n��{^y�¯������у>����2��Kc��=[*�U�ù��(��K��.��M�A�ĥT�o�!.`��o'�Y�B�AqK��F�q�����K\\�c���dSL��>�oTЦ
�F�4�5]b5'���g�rN��������N��j�t`���B�@)#��? [@��f�w P�Ok��v�Tn��|��"
"N�Sx��w�++��ǧ�,2��7n�cB���X3�xzzzvr�/�b>�?{����DT<}����TIr����\8g����1��� �x<�Mg ���|�=Ƒ��׽�<8<81� !Fk�n$�[ �:0_�:��:�u-��!�U5�Ά���`PUU�x"CdWTuUU0���R�YU� 2�"1;���� ,�W���)�xA�(Y�TRfy��Oe�O\k����%�.�����8�y-?���s����yi��t{��*��b9��A���Ѣ�����ҁ�ȱ���|. ��Ї���bLB	鯜-'��\��	!y�R�~�n�U�t�|\�@ �v,ӡ>��宀 �e� [2t�J%��k������x�4����#�$Ҷ�@K.�9�!�N���Ak?ޝ��S!bQ�}#"UU�u��Eq�yDd��1�P��t6]Y]A������-/��W*6�����td]��"��Bx�f�t Լ��F�W"�b�Ǫ�ff�ܙюn�9��> :犲��9��̫���9���FTߐE��	R1#��bXc��I�>�(�% ��������JY�  Vuu||�����t���	>h  �H�э�}p�FR�+֝���_�O�����@K��\�9\ �.}��:��[��B��8�&!`�J8cА�3�n#v���A 4A�!u]װkvnU@�3i�� ��,��.�O^:2���M�$�6Q1u��l�����T�I�}y9�_�%ۭO�C��(��7��Ej/�-N�%˵���[z\h/=�y�-��ރ������tYT���JW�Bf6D�Y����Ǩ3���@�,v�,��$�-��"���qy��L��VL�ek$/�4���O��ߵ�� �����o����}�ޗ��^Ofӭ����o�������= p�E��\��X���������{��}������ַ������{�������w&�Ƀ�֭[�y|v6���V���ק����������כ�O�����������g�A8�.��Ul�sH��u��H҆��t<>�V��a�?  fv�	��mХ�*��c� ����3sa"�D�����O{\��F]�;3Y�Nk���.����v��(�=����9��8�w%�3�(b��B6��`f�x"���y��6LR�?
j�Mc-��(���ف���i�Kd��	���XKZY�x���W���W-%���i�:o�;‹!E�j�q--\�\p���`���I�g�qP�|����j=p��R\�u�w�QJ>�� K�k��ːQ�'@��Ґ��eT�#�@(MQ!c� ȑG������l�ݥ��K�Tm�BB��	``��X�[Gw�����΃��|l�,�Xn,����h�}��B��˲�+
���4�����"�ɤ�+�%��Ҟ��Tx[D )�`�p0��z��jA�A�[YY��Ύ''GϞ���u�"��C ��K�恾Ä�\6%RXBZW�8`�PMBj����
"�6�J���� ��3 8�x��K�e3�H�2��9�$�sJr��~�(,͍���1F����5��Ө��\ᬳ1�s���Y�Z���Zu�>�٘v����[�b�]%}�s��=�ָt�I��  �."I����|2u}�<+u��+�B�)�;��V���u%e�s��[j��AuP��$�r���#��ZFkE���NUu$�PC�Xj?����2�N@*�"���I�R��l@cd�"��) D���s��k��0���3��Wou�c4��݁��""�N�j��	��d�QI)'''?���N��{�zo}}��k�+C�s�j:���_�������|p��[~��'�|��;����O���O>~��7����8x���߸�ڟ��޻w�g?�9����?n���>��|�;����'�����{�����������޽���~�������?~��E�X�z>-�m�LAB�Ӆp(F���L��iF����y=�{�~�_j�i�����+@&$��wCdT��P���!DAM���~)��s�?�޳��X� �*��	t�]v~�^��Y��y}�#�&������pZ��!��i��JtG�\��z1�J��A�.���� iUwn�� �}]�?�=Y"��1�:|�sc�����1f_D�]

 �ןs&1�1�a꠰����ِ��p��޾>���!Y��wזZ�R��}ڤ��@&Iy_>�ӡ۔�Zݬ|E�QkBR缔��T*���bE8
��Lf�Ѩ���_�H�iЎ�$ٖLW�T��� ��1C�,�9rf, !�`���0�Z}�Yj+e Pb\��64}��t6S��vPr.BDB���pr\���X[�`8U��^��Y��EX�"��1��� �4�5m�rd��1A��w�4sQ���	c��c]Շ���g',�9c,1�Df�g���w
�*u���k�!��$��.o*I'/�b-nJ����Gj�5\7 �� R�$!z�,q��*��"���u�E��l>+ʢ��j^MVWכ&��; ��iLX�6�I�E˕ʣ��I��#w!  M)�E�X�������Ig"H��DW,NR]`&�_�����;w�h��7._3Mp�q�n|��՟k/���w6脐�}N̆����EL��}�>����C��Cb�E%�t2�̑�E溮� �4�9�0HҮ��pa�$A��NS�-�@LJ�����\�hQ-L֦��h�!�	1��ｆ^O�>�}���ht}��������_�/��p�:������pU��Z���=����k;7n����:��_�~��7�X][���z�7������d:]]]�ns0x�oݺ�����~�_}�a�߻}�����X����_���d�o��,#s��y~��U����lH�Мu�52�� ���9*9�D$bV54J� $i�f{"b�V���y���j�����֎tWb�!-���N��W����(\%�Թ��S��ȣw� �dCZ蠳Q�A�p �C�J��� �5�ȍ1@�H�b�� �=˿�C�H@@Bl��/�@���0�,��G�m�H��DfQ�TH2�<TU	%2�D�Y �v�j���  �V_�y" ̂�Ϋ��u��������.<��=��Wi�o�w���'�>D"
!�ש(�z
�1��j�
���R�zwv�u��iJ#��.�ȑcD"C֐H������N(
���'CD,��Z�̚؍Yh�l�He�E ���>::2֮��Ƙx0�����3�Iɕ9�6"$�1ӌ� 3[$QҀ�s��Jk� ��2eY���c�L���$�dp���J%Bʢr7��<k�@[�����  cTskse;���P���0�Niۈc��)#�)�a��_�
��9'�ƚV�9�QVT��s��"CT8W8�:� [��%�q�yc����ne�6��T�H��@;UiZL�*�8~�$P�|D���s�����i/1��ۡ�"���V~5u�wʝ�7�����^�B}��S۹98Ijl��  ��脴��(��(��i��땽r��z�ee�O"�)���G�fA�e�@�0+A"X�X�LH����,`����"�M�?��`4\_]�����O�������֚��>��ۛL'�a��������/�d���������x�/���������j��o���u�?z����?>>>�1�������lnn�>}������3Dl�A�ԥ9&�����ⰼ�h���� N���l>��E�1F���H��;�&�T�9�DV� hUl����9�
�w�۽S�p�u$��a������`�n������������;�g�Ũߥr�6zc��e�CK�1�8�|$�!wc�׌C�9*K_׋e��"_!��;b��>��m�J�w��%�I�2N $C�F3�&�h[�J����ӎ��yM]G$Yy�E��5���55S&%`s����m)F-���x��e�y R�m�bp�X1nDU�1��u̬�D�%�8?=�16M��S6��"��X�})��J�l�����,MAba����(]�P����O~|;&m�a�3�J�l�D$� \�W$ 
�!F�u�4���11Dk�`0���u��H����X�����-#	s ͚"b�j	�:�e�3��Ȇ����J�'4ٟ`Ba	̂Qb�ER큺r&!�����pLmJg~��Yk��&�1�S�:�bE�|L CX���t�B��������JK[=��)̂�!D1흆  �L����!��� q6�q¥@	��4Z���_N� �
�.���"]�,�RF`֘�;�D��s0��6�kUDt�^�t�������Eyoƌ����.��'�϶9��&��{g�[�.�yᾋ�ڟ�4�����Zt�[u���C�7��)��s�(������ØM�0�JΪu�����Z_��n�Ӗ�q���vJ.(S��"�Q��fv�1Dc���PRS�1��O�z~���G����vv���zea6����_���1������M�C�<���!́��Ǐ�ſ���2�NC��G?Bĺ���������7O�<A��~������	<~t����Y�5Zԕ:^�#�9��V%�IҰk퓎�^7N�f��dH��ON���~Y!��}vL���#+Q}�(���&��H�[x	��e~�eq]����aW_�%����������BfVŶ�*
���Xs�o��v01��e')�4�����{"�ʋ�c8]1K���1c�u��S� ��o�a�Z�K���X����X�W�f��n��*"&7�ц:�y#<�"�3�U-�� �G�VjD@"醔��� 5�V��Hg�P��I��ڹ��R���[����Ak- ��^�+����n�3��d�U]"��-z��B)���{,�J_��1�(1�#���!t�H�Db�E""�1�gm����$yB�"/y?�	�����8k&6��:��p� ���ʃ0�y5�ͭ�h:爬híTJ��ֆ~ɛ�1ZUe�!@���RE�u��qC�ԩ^0��} `��,QDP��S������N�4!)��[���怢��1b��.�3'qQe��,H����� >2!�r�6M7����D�|ӬY��:������s��*�07�0��&�W��Z���`8\[[;;;�����yU9k+� B�2�(�xN�8f�*�1T�@' (�� ��\����l�� ��J1�֓�o .�_���!�]��N'�o�՗��ijvʶ�""�d/�T��qMh/qŁKsDxy�q�Mՙ��`ee�����p8T}m��. �dqd(���p8R�t�M�%H}�#E����Q.yv=����@�,��R�lZŉ��������������/���w�ӟ~�Ž[�n}�H�b{�{f��d||r$�~o6����R�+�y���C�� ��DT:~��n��j��>�S�������h�E��S5VL�"��k�
PI����Yi59��ޜL�>4��!��x����9�#`d1�Q��L�̙u��W�$��0	�/%�A$�W_����ם9���/N���aδ��?�t�^��������`���]悉 ��P�A`�01�o�+X$�@2�*���GJ�.�`��U.���(��Sh�*Q�nC�%4�
G��m�ʕGwx.�,t�9D<7�4_�@K1��GB���V_�T����^Ű(����il�|�|�{H�����k�p1��Q��9�� ��O��Faf!�!��]��)��uNS�e�G�G�f Z΀�P!E��(�r8�e�/�B�Q�:Dz�T�k���̪��r�5��1����އ"!�mD7ccl�W�v�&"AR1L��wI�q�ξ:xn��"����6���6��뺮��`�R�����P��h $��r��B��آAE4�����nQc�yLh���� �2Ӗ�El1�e�Q_�(Ĥ4&@Fu�6�y�	n-��	��n��};���s
V����~�k��>d檪$i8����
QD�uu6W� �FD������XDf��$M1�,|�A���"�4��.L;g@R��tc��t|A]�bЈ��~Q���ކfC:7s��vᕋ%��,���'����n�Ō"]ed�_���Bk�s�Ҙֺ�"^�}���3��d�y��$e�E�]ubI�uu||��lUU ���D�Z�Hq:�?y�t|6aW8D�N����[p�v���HV,"$^�6-�c��v������о����)B���ib]/_~��Ç`>����?��L���d��	LH���8��i2Zפ善�κhc��	ʲY�+Ġ��4��*QQ����a�������uO���:`���
�ȆP�8r���g]�e�y f�>���S�{9g�����@hE`����jPK/|��ŗ֟�+��$,� ��Xj��d� ٘�*�dU������1y�t�s��fz0���{�="
�n�Yw8w�=���gYb����Z�������F-"��`��,�.�+�鈏:v �}��q�Uׅ�u��*��}w�PF�K�ü�������``��a�O;ח=����i=
�mZ&>::z��q�1�U��ˉ�Z'5{K��\�N�[[[��>�4�δDl�fN�%��6���:���P���S��W���©$��!�5M��=,i�%�Z��"���8e:T��ߠ	�'4��hX�o�)C�q�S�F�C�d�X  �%�V�
8�&g:�lEӶ}�w]g
2�[\��*��+rJ�&0�<�ں���\.cJ>�O�9�&�x4�㞙����D�R�Ѐ�D�1�P���@�ͩ��wJ@���v#i͒��� �٩&*<���S�x2iK� DcRD�B�	M�́	=�����=�/e�tw�A<;�K�cQ!�[w$����Ѩ'�m�!��/:Q�Ȭ�rC�(Vp�Q5��������>G%Kw-����"f۹;@��&������O���"EY,�锉'������i�J�f�n:����OOO<|4�L�v�_~��!wdv�p�Ů�Ƈ��ɦcA�ve�'��{�
�K��<<�-gQe�H
%΃�I�S-�Y���;j��\���FW"P��~�Y���c�P�J������Õ��Z�z�X����:��q�ضF���:�w F��As�~��߽�qJ2�/���t:ۚ�v���=��L!��t�����?��f���a&@���́�/Z}"u�R���D�&�Tϲ���Sjd�&���\�p�u\S,a#�5��o`MΖ����Ҁ��r�B&@U5�hm�FE���J,"�6- t}�ܶmMcʒۦ�Rk\mb5bёx^K�H(�	LT_־n	Ld���S 㦁���ĩVo� F�u�2Sձd{��\�Z�W�繞g����6IL`Db�i�5\�D�'�Z^��D4+�C@�kZ��K�.���w�6 �ﰾ�=F���D���]��]zz�\-SL}ߵ��t2��Y�Ҝmr��?��ݸqcgw��ݻ}�7m�v���a�s��H��s����tl�ﲴd��#�a��؋fu�qt�ZD�E3(�ϖ$�ι�+y���Ӡ�8	ɚ{T#RQiP&���'t�^k�Z,.����\��Y�������OC������G����{9���y�LJ��{^���)��ir�w�|xzrrxp�꺣'���r�;e"�L�Kj^�e���E	�BPT��ì*�&��(,Z��RHDD鰊@���"��+�F�Z��S[��j\ׂTL^��HV"0 ����`!N����8pB��~Y��@2{� �
H��B�Q$g(��6�"����1#(y"�h�۟!���N���6�O2�rfb�AY^�qo[+��t��&���P�  ilc��pmo/�4Msppppxh��HHV��}�Ȗ�����O?�1Zo"m'��c�����^O�0;hAۂ�]x@D�^O��8X8r=��J�U��~0PT%�rEP�R���
�N�X�
�
⋞<Q^�RkeG�B��&�6����n���Ds^e��F-�V�YƎ�Č����UQ-l~�5YG�h��b>��1 � �󴝾��K���{���#O�S ��ާ?��{��ܼ����Yk\ǳ��S������U�)�gޘ|D��j�`���ѻzl�l��Ng��봔����X/ ��B���;B��RQ��oچ���[�P�y(��?s����� %̬ QM)��*!a@S���}p۶�7�d2��V��bM���籈j(�����4�RZ��"}�4~�_�2�NHƌ���p��������u�3�B�`�B=��0��\L��)כ2y��
������ѣG&�b�]����}�ۻ��Y�O�fEZ_��i@u�X<|����$����bJ��l�$���>�[�M�p���^ J��t������/V|p�.JT4��R.̇��8���BJ։����f���*Z�*�/��;Y��BVta_���	�.�l��e�LgN�V0��U:9>>::���]7��SN׮�߸q�i�v2c�!��Ha��r9��sΟ|�ɏ���	�층5-;ݬ�����J��!�XrM�0�H͉��%�ضPP�1JήBm��;�����1���+��Â*v��7��ҍ��N�퇪p���\�U�d�_�##�{� ֑"��
���-��)��T-�8���W�� B�Z�o(�)�<b��d"b�[�lOy�j�^����	T�|xVO#�0�)����!,�2�ϭ9";ɾ�M�a׭BRz�Q��bD45iK�&I���s��N%� ���m URKk���d�Z!TBFbʣD{�9Y"�jVp�,0��&Q9@E&���͙/���"��ի
"J�nG��rè
�q�v5l�	 �TP����6
�'7` �V����\W�$��� Vڅ�EE��L���;e������	��xYMXA@K�L9��l2A���8��h����bT��^Lyj�T��b�<21=�Rdǳ4$T	GQ���d&V��hn���c��K\�,V���֯ʍ�8J�k����3�Z?P��;,�"�Yi��L��+����5�%�H&�l�k� J�t�ꇲ`��)*I%Yu�֓\�BOjŮIJPc�֢U���ߊ]i?A@BR��.�4��O�ɠe1j�)��y�H(@5��r�^kV�'�<���m� �4�m��lvppp�����-@L9[���^ ��1�����u_5�U �#E�R��5��FϜ��Lin�!I `NT�r&2<�h���i|�DR�G*� ���e<?�"9{f^I�����Q�2�v׼b	1�s�֡j\_Rd�bmp�����u��aigP�q��qWĮ�\n�^�eOD?�0A�dM�,�R�̤J��e.����ׯ_�1�bhB�'%�Ӷ��r)"��t��E�&خ�n�k~�͎!�<�_���۶E�>�1%D`fRȒT���B��Mf8��ힰ�N؄ 
�@�9gz �8��\�V#{�ܩ)*��d�|��$�a����D �
�\�TߦŚqId��C�c��Н˵��c��Ƿ�O�}��s�VU���|ZU)�qx�iB=Q@�ih���W�3'����L@\�*��gggGGG�YQ��d
9F3]������t]�`�4�Ŗ(���k+V-����>�V}�8��qfz�;+"U�KU�B�� ���� �`��R$�"y�X̻.�4�N�����ൔ-^W�l��A�4���0�n�Q�/s�e��+��aU_)���	��ґk���rrr|v~��*��<� h��"W`bsAEՊ�,���]�0��5��-D�f��?��bS��]�D�"�������S8�>/*��C>�SJYr�0�Ѿ8@I����pkaS�����1��.5�Be��5Z9�Q��ku���x�1��6-sh� "1���A$#ځ��a�@��������A��vq�K<�yͬg^��/:��8�f<Y�R�/W~���5�
c��kX�
�� [%M\.���3��Ō�Rb��p��|�>4M��J|H6Zi�;O�Vc�J˷�|^�iƽ%M^�`����
��ip�#�.�][��L�ư��Q���"Q$�Fr2��ʺy'Y �
ͨdi�E�\�������*z�G�DdE��Q
�&�j+U �t���@�=C��5�dti!01s`R�`n��a��j��񣮋�L�L sV����1ƾ�Ch&"�n��Q�ӞA�Y-r��h���vt���b��yƲ	�T%4��g��i"-�؈PD2"�^.@�q��ݥ-�'�<�P�fE���q ��3}T՚Q{"o۶!%cc9��͂.N������k&L΢e��u=V@P����>0���mLrW��wd��ՁD@�?MQUc�.�*���2enz�j	����Պs���3�Z�'3��mh!��TN�O'��̡i�������8ǒ��@ 26��W�G,�@3�*�U�XwQͱW�v��@e�1�d�Ո��E����"`�X�&Wr a�`��
W}D�x4�ӍGr�6X�W�M�X���o�p��vlֽ��_��jD��uQ
��+x:��PF��T߼�^�:00���{����V��e�<�ci:
c.�j.�%���Ȥ�JR�7�%�N"S��E��M����T�+S�޼eьUa*}�K���bu2]����XtF6�~E��ڶ%®[�"3��DUt�qn��f��YT	Da���y�ck��0&��n����iJ����7��>l��C�5�iQ9d�F�WS5"�0�Y-VM]��5~���*�������ʊ)@���*dɠ֓]�x:���k�D��'���hb6���?_\�#F��ZD�Ŭ�XUd�x�U;@T2J�:*�A/��kK�� Q��2� ��-(Z��[+8���-���\6q���6�d2	M��z��K��Y�C"Q"��03�.�zT����z�\�U�>��0K��(KUs0S���ȓ�'Rڡ�" ��<����A?��А�Lp6PKϽxF.Y�b�30 X��!�KipZv��!�`�w`D7�#�b�f��E��`���f��i|��Vr����|82�L�"�ۯhL��T5��ND�/�YO!�6p���'�Z"[Z���e���C�VV짺��q���U�B&��~ϑ��SF7"$�k-��M,6�%�"y�x�rZ#���"-�	��6!��G�v:��U5��mSJ}!�ZD�	ER�D��SJ9F ඩ�Aϴ�*�g�CDD�ډ*������|q�N���	s�5��̥E������6'+���H�u)%�eP$P@^-��^r�TAI�Ƹ]+���Sht�5-�XV�鳴��pY:��g�JsH��i�!Y��7N 3�!s�Zf]�sU`�t��/^|�^���%3`���PP*�:4D�x�a8c��2l�f*�9�&4�A����Ъ��-���>�'��K��i�zy�1 -���2�nU�����5�3c\ChBӨ����ӓ�����^m������I5�>�2�2i��R �T�X��r�K�+���kmzG�U�hީ��5�^K�v�zzF;9.P�z�h
j�KkrT���u����C�jh��]U5�K����O���A=�rl�^y�,a-�G�MIRӂ	/�b*�d�:<
��[Iӥ�%��(��u��23�v��*>�ㅐ,��mB`d����Ϫ�j�
�k#DP+Y"��ZA�E���9���	BMhL��cT$l��V�T�5�J)gL�$Y���w���;>8��A`$�v��b�6��B؂oߡ�ǂJ�L��ڶ�-sFCb��3�
Q`V)���C��"��ΒU5`������T��KE[&ٚM����vq���<���y�{���xy�݂,���,T�H����^�ơJ�!�����@8i'�i�%D-�@�M��Įͼ ���C-.�ΔEa�8���u����i��e�aF�E���'Ѭk�?R�q������\��? ��	��	�E%�ld�V��Y���@����V��\m朌����D�il��vaE�.��*u_>[+9��`�p����ɤ%bu�E�X0�H	'mK�n��k�j�i:�2{ �ĬY�K&To�� $%����Zl�Vs0������Ћ�c�e���R�#�6��-A -U=k�`�<XK�@��k�K��t�{��g@2�V�blu�^n
��-[��3>��� #�:�v�ڤ�'/፺�t����ƾz婩��Tc��Xa��2�)�>�n���裶��QD2�5H��A�iS��8�&Yc�$�S�!p�L�������|~.*�g'��DwN��$ƺC��u������w�C���5h �K��6�~��xJ�װ�7��YIe��F� P��DU��������QF@��ϼ��҄��Dd6�ƺ� x_�XE#��v1a,:��\Ǟ�u��1Cř�������I��*�����F�𝨪x��x��	��wmg(h��4Q#$�\;_����ş�-9��k��5���) BV���^��#�$)+����lݩ3�5,p`PU�jg�.f�1�krB	�}���ϴC8e � C`"��C�%�d ���̾�I"3S��hg=K�14�"!phB���i&Uܥ��2p�1'QRfVP�}	 
�D�ɴ	�-Nղ��J�TUP##��p4a}#�#����zg�n�Aؚmf �&b��<Ζ��r̍�k@�0k�"I��H�	���q���8��J���XlT�E����e{��GѤ�/�^��$�)eVE TR�p�����d�R&" ���kN^,J��f�1�����b���k��
��b��^`��ܵ��J\� �Y�a��^d��m�Vu`��V���٣�{���က�	�$Ɩ��D�����xbm���N��R��TPB�Ev��x`���EFr��~�2ߢȱ�Y �b�"]TfO�ͫ�\�P> �`{�?(�S��n����IN�8HuT�[��{�d�Δ��J�����U��Z��b���Z5Ӧk���"(J��=�i2���4����﫧�C���I�>��X	fhS~;�ͤm��{�U�������m۶mc��md�CQf�JLIr�ZL�� �r<�k����V�3~}�Ʋɜ�@%NT���ň�>E����Ðp��Q�Ru���l�(���zXYk��X��@i�áF�K<������F�5u����C�b$ �
�>"�&�`�C�b���jb^�Y]�k�����,�,�Fl��G�Y7p����f�gM+�PCe���k�K����ɋ��Y3KE�9���GT򯒴
]ߍ��UI�Ec�P@0nHK4T�P�T��Q�mZ$��#�{�F�⮸.(P�T��!�*2P���Ql/�lHI���V;u)�m�1üGxYYI P�O}�u�����,�`�	e�;գA$ĨZi��мk��$T%��Ғ������ؐ�2�(03+@�)�h�}M�#B!�p �~7�`������V�	��d�}
`�йBy=7�B�A\yԇ�u��
��v,�7�����Ջ��{�jU�������9(Xi�3EꍆmHڶ������M��	�oa�D�� "�D���x#&�w!�<A!����YA	�f�tBJH�՝���C ��M����	Q�S��	]SQ(��gF��EQ����Kf�e���z��Ѩ�=�7�J�u��W�ٹ(�+in�^UY@�JT�p�
8����R���2���T���]�Ǯ���,b�wU�Vj?~(S*8��XYHu�a,��#q9B�}C%�����Gv���+���/Dx��6Y�2`����j��d�1�V+D��f"zvv�����/����c��� B��5? x6k����͂�:�h.����lW�]-Ѫ}�<�o��,�s���/�g�����4�%�P3"��~'0&��!٤�oxU�\5d���En��p��`�#j�����oe��LM�e����!�j0_}��j�Q�ڶ�Bd�A���0���E��ŧ]��%﫨��A�48#
R�>���)/Z��e}, �t��ó�N��d&Фd�d>-&��$����z{�j�l�"gs�����f��{iBpKλ6�b�ämo\�i�GhMqʮv~)�T?b5���� b(MΞj�+a��О5�"�&�@G"��1iF�!�	K��Ѻ��6�`���ӽ����5��>����_��K�:*�D�Z�`�2츑���q��� ��3��'�h���;1��I��mfR��
"P`s;��
�=�Y�1�Zk{c�A�h�y��Y<?ǂ�P���N �൮Z�5 
��=�P`֬0�͍-ᇣX'�����(EE ���2ڪ������_��C�t4
-m��=-,��QZ�\ l���CY�U�*S���= ��%KҔcjCf�V�X�˖�<�3�B Ȓm�)��-�W����)r�	.�EpH rz0�#���q�n6-��e��f'�>P�6�W\�}T��"@���.U]mCW��ҷZ��R!�᧘��FDk-c
����Tv䥌�5��ylnS� �(:��R�7����ID<�������ۗZ@���f�����*�"��-�#�n������"dl�d��P���2���Bh��YNi�X�� �mڜ�뎎���������/^�JJ���m�9�lE����p�2�����~(����e3^�:��?Ѳ@�>�f%����u��
w��{hm[Gk|W6�"�:uj�SqX��G�& 9Sa�BT,��	I�"��E��A���XAK��Z_�QE��w�jL�n1�Rz{��"��vT�b�tf���4P�9��(ύVmrջV���)ʹ��b9U�n[�ܵW8���úU�t�����動KT\Σ�#��`�Z	���9�RL�d�,"�v�ГR��Yol���^3�h�@����A@��E� 7�lm��FG���ppm�@ =�C4�P�9�������lE�$E����iVFp�NB6�΀��Ř�RJ�G�:� ����[������=�b��=��9�K�݆^O�aǰK�Fϼ,�	$(�q�� ,X7B�}k�m�����P���b�E,��]�b��B���Ch�Rs�:����q)`���
�V]�{.�Oq���o�6lDdbOܭ�Y������-\�f�\
ޤIbN�r�����Bh��P`RJIACM�'�Kb�
@�s�}��&X��������o�����EW� 
h���%�P���@5ʾ��7�BE��e�w�[l��^0Ьn���s]�ɥC���03���4��*6e�Z�ɩ�*^GSྸ�8��� ��R0�ŁW��!�0��`t"S�HU0��f`�.��/����P�aБ0�h�mjY���7"���"�Em١��^�=�M�J��Nѝ"ڶ����&4M3�m����G�N���Z���9�Z4���������oO�S$�؛�Y,%���||���Xԡ��<�1`��6t��z�'�Z"��gU�
�8x`f�W��!:���\��ܚ�D�T�vo�ƔEDC ���( ���J�43F��	�E�j(�f��?:ޮ'���@R��J	�p��G�a!5oP��RD����8��Oķ+x����e�]� 1y���_b�v�Y/���m���#/����_PɊ�@�H�lȀF���E��{�����b6! [E�5�b
�,FE�m	��z'Zo�D��EJhKU��aS5!4���a�����WM�D8����H@E��iZ��u�fZ,�{':������ؗK DD����E�$��E_�H�L��ʒXGk"(��B!�*n � 4r�-�,R�:��7�a��|4{�3��;;rD,�%��m s����5p-�(*��f�^Wi�Ή|F�n�����4�����ߔ�D����iP�x���e�J�)�(5x�C�ˍ[�U�
�"�%��є��	�������~r��NB��H�n�ƣa1j7�(�g E����o���;�L�Ss x@��� ���Gw>����G6�}�qVu�^��-�M�jcO��61e�"!�|#�!�&H����b̍�3V~�Jh!��xUq��/`wUN������=�ȵ�j��=G�C0B��S�D����.�x��;k����<�����R��+fBU5� �l6%������B0*,C�/З�gD�fj��5G۵�:�Z��p����S��F�
#f������f�J}Q[�gɁ{E ��b�ä )��SMA$�tb�to]�V�''����l{{��\b���ե�y }tn)�TY��5�x�/�I�N��+��8��ݬ��d��H�{�CƂ� !8�@�V��6 �r顒�e*�RV}EV���_�T1W �fQ�%��i}Q]	2T[�~*�j��"8��)�2f+3�t8��!��pks�{�ҽtե��E}��բHMx^Tak/��Cņ�ֽ;���a��b�_}��#!�K#P�u�7����f�"�R�NH6	��b��)������,��E�;�)'�و���MU.��22�d*����V��As:�Uck��@9��q��$DA&��p$�.#g��`4���H)֋� u��ά�vl6=�e��Z����ʡ,��a�e)z&�&XR�Vꞑ���L�ID+��G�68h�����I��1F��&+W��!�!Mڦm�(eC*�/��8�eb�\$�T�W���AF�M��V��jB����l�іP��HZ�Ѧ YbL�FX9�8@�k����׶���^u��"tS+�u�_(��\�kY��" 7!��޵k���_���߸��GGG�sBhΪ�U����B��'��s
!a����,MBU��JE'16M#,)���s��!���r�f/����� ..�ח_��#����9'��WQ�D��Ë�@����|�t�OAi�1����RM�Nyo�}�/F�Hؘ1d���-;��7@P��X�2Xe�k@,A�"���͛��ů0��������J���=��h��OX�zv9�5�	AP4k�a�+֗#�L��I��)�2"5����7�������poo�[u��M����
��db��'�aju][�wD-�����8b��t҄ƕ�(Řnz����t���&�=,��>�*�E�Y`s�,�d_��Ҧ$�FC���A�<���V'՟ӜU5f4A*��p)�Zz���B`F��\"u�y؆�~@�brz���s�esx��4~e��@A �Τ"�䃃�����y啗��ϗ�ea�\ڂ������S$軮m��l���G��x��)X�mbB���̲1Z�#{1��dM�q�p��13�JL�zo���ۦ�Ե�O���.��i6-����V�c���:**����>6�X��2�؀������%a�����Zb��� Z����ɥ��:VUk�9�ͺ�)��<���H�5[�T"S(0�k�� �r%!'�,�Q봠k��"T"0oC$�@A'V���38h�9�z��6��2j�PM�-�bds�cG�!	T�$�I������|#K�Cy�%$�(k� ~��J�q�z�z ���r��8��Ke��2϶�����;��x��q۶6{e���X�b�9��-<��� h�	T���9申��ҏCh+],�(��dQB��%؎s� {HQ ��� ŇDPd��R�|��z]�g|w����-K�����! �+Ѳ�{� �Գ�K�T�VK:J��S�r�MV��V��$����77��э$#��:��pu�gÈ���.F)��Hؿk�����$�z�n��-!#7��$&��D�,��R\j5!��0&�$[)'L&��� �J����>?ۚ�����������f۳n�4�Q��l֘E1�d1|���a���kn�Z����ՔS3�T��s/9A�
!��iJ�V�U
`�V]e�Վ;֞������Q߲�2U���4  T�+W�e�K�� OB-TG�:^���G�P7��"��nT�"�"�g|�{~����7��]����ɇ_dlV�@�xm�ڍן<y��{�V��m��W�2gG�T$�hM���^=88�������� `ʹL��H!*]��CdI89K&t�zf^����쮔�,1�U�"���M�U��x��P�Z�A�@�W�����k����9�b�����l�-fd_���6+'���Qa���B є���%��d"�aW��hIEs��f� �T���(3�݁��i��X2J	�x
r@�涩���Il	�.�`|��Y��'|`�dɥi�b��2�T\LUk?������{ό(��>�&8�mZ���-(F*k4+���``��� FBԜ�Ԛ��^c� *}�c�a�53^ �cDo � ^D�"yT=gx ����2D��a ���J�G��;�}���_|����I�6�<i�ж��[6J��uJ�npVZb⚙�}��V�5�V-�R�9�5K�������������b�4���d�{�h�V�
��F����D��<��R�L%�̍[���T`D���/"����wGd��@�����.5���<���Ɔ��c#���-��>3}�[V��D��B�@vV?ڀ l;��3�L&�9Q���K9�*Yi������%������0s��p`"f�B�JD���2C�"�f:��j�QU�ݟ�jVȚ�.Ǹ���=����Z��J���̈\H
�-G�����u��L�UsP���,`n
D��u���D)\�Aףȩw�(%}4�
b ff��Vk�%eUoEkݥ\ ��	͘=�)�����~|l�g 9����.�F��w�	�լ���J,A����v�ⱍ<*)+���R�,B��ƅ�ui�UUZ(lf�^>�e�Yr�Y��-���?�˿�KB
!x��"z�@�����������{�����"b�Y���9`#9�}�%3���HZ�X�+6������	M�PRq����`�%�ZRω�-�
KU]�~*�1�M��&qU�ܛ��L*@�%�("l)ԣ��:�:F�X)�jz1W���iu�*�N����Sg<.�s�`�&� R�^�� `1���mK�?��DH1PM��x��*� !��1´� �{A�s<v`��J�$�Н�(��*��Fu3Zg���ĂkO2�'|l[�%� �8�ʬ�+�ӂ�&^C�E�vU*���БtN)Tat���)礪�7n�Ȓs��bqrrb�T$&6�~�F���c<D[�ۓ�$�DDmۊH���8�W`P��U���A$��O���g�n�d%:%)�
MhVE#)d���G�bT�$���-��ܤ�5U��Ӫ����=������D�Z���בyIc��QD��9���>���.P0�S�.0�|�rrp��v���_�u�Ϡ.X��ů�*�{��r��Fy�+�5Ir��Qz��7�iC�,��{˂bZ�R*Fc����a*�p1c����mc{��)Sfڴ�>�����`�����^���$��Ų�$�3s�4��u]�qT���%-@����I��'mk6h����K��EPE4e�@Fg�,\��7/�� �N�#���)gP!�m�m}�0Z�U4�%��
�RL\4M����>�|V���b�j]}�0-Xi1�ٜ�g��V4}x�2K�������R�/.���!�]ū}�K/���ō{m�y! ZO6��Ѯ��uE��M�S��3���&�	�`6�s��V�ҭz�҄&�d7*ST����/&��|a��Zbw�{�zff�m�!c��~*6��W�5D��̓�ef��ú1FjGJ\�O�X O����c3KBr`��	��I!�+��߷�b�9�0,�;?P�WB#���8��?���z���uaQA`朳�" �fc�B4yŒ�T� ����ҨD�����I4���LA���l�)[ֶ�(��wվ*���!4�	�4��Fd�tŰU���u� jL�ؠ�u����-���1��p�BKCA5~�"U�6V_۱����Ë�Lղ���F�ģ�  #����|�w~��������O��}��I�iҶ
0i[H^F�o�L)�����K�''������u~~����dy���/W�c���(��s@l��qz<���$k��� ���"���D�l�GɶuN�&��eW:ɔW�y�uf���{_��>�J���yCD� HȖv]L�R��|�*����Et\��t�r�>3Ƈ�ϋ�]]qK�[�Z�}E��%����Q����:��^��T�q$�3c*ů�lw�0�衺v�R l����6C��*
���±��@�[������`�3��ϛ�f�P���5P������?Nu0���Ҧi'� ̉�~��
��?>>��f;;;׮�goK�(^���/,``̇U��XڠO��RȒ�zn!�r���@�H`j�4�Ų� E͞�dpF��a���R��,�'dK�P���R�JT ��[S�!f��%L��f꘳~x�:[U�+�Ŭ�8-#|Σ�i���n8��Z���-�ɜK�F�陦���t�ٽq=�t�+�j�Z���d��d21�a�N��ӄ���U5����_�*m϶%���/mmo��h?e(�W����۶m�@D��1s�s&�q�#�"���@1�D@��;�L��0t{*�e�%E�����n�I��A����5�u��k�F�Z�4�I�e9��u�*(���~���h-�U�<��y��Ja1 :�񄫪�#�0Ƽ����%�( ��C �%,��3if" 2���%Ricr	q5��Y�*2l�ٛ�hq�,�6��y�-�f��2�j��BQ��7ɉ��fw�+`�^�؜e�k�E�h�fDH5;Ҷxe��௻\@!�}|r�JP{2���d2 �V)&?��Y�?z�/��G��<�LC/ "@���y���YD�Mۤ�fp�J��Zs�Zl�$1sh�r�L95m�pӶ�AZ!�a0 ���z��䔄�Q!4s����}��>�� �f&62��B��!"Y���4ޠ��Zĉ�D���i�Y������ui�(Kz��.��bu3wF��J�Қ��3��"��X6�"��R�Ѫj��˫�
т/�v䔑�q��"DJ���fh�h:d�g��v(�����.�Ra����� �"c���͵�訳Ș�E�Ū�䷟-vmIo/�*�B9瘒����b��o<@�fJ������t]�S�cT�$�e���!s� 9��"7�.�x��%�r�4%�1��?	���:�V?ߎHd&B��KB@ť�\u7+�x&��=�́��90s`$q~��d|�NV0�_ �R��� �u��ڠ8��t�q�vu Z��iq�ұ����>G[׹��l�g]�Gg� �f�k��ĺ[����C�AbJi�\]�~�����~��w 5����eխ�- ������·5�+�c��>��BYflS�4.:�y�u)�i(
��`cAhu�n��ڸ�Ci�*V����0b�L$@ͮ�MN�%bCE7]��_ʮ���xB�!X!���ʖ2�4����z-�u� #>W0\Q%K��H�4A6l�z+|��Uud�ֽ�m���H=3[�g����)*wU(j{$��7,J@�(��d?��_���D@�Z�%�R�\sW�dq.Ԛ�e������a�-���:�-��l�K�s�VG��q"�=��I�:5E��	<_D=�IEd>�����] mے��FH)��	�R���&V��4M۶]׭V���Sp�� ��S��U�(��GE5!P4��ܙ��!�!���)㭭�$)ƨ�HD���$�hk�LB��r?��ts��-�����i��&�N��y���w�'�I�ꏎ�>|�w��21 �C�ɷ������8֙�K$3"��KW��������kʅ��md-�j������֓izԕM�P�j	<���mL�!ƾ�{�،�u�������3eײ�8Ť�D�;kDJ*"I���ʈ�b24"X�x!��*��hW;�A��g�Xl2<��~k#St8��O�,�����]tj����X�#d	��fg Y$�Ehs��i&�Iι�z;)��z�v�"�|��rN�n�U'�NR�bB�\�Z_��$�J7���Q�zd��z{l�v2� Bʑ�9����y}*cB��0B!�dd�ƃ'T8��8�$j��U�iN ��B@�J���R�����̜�g,�5
�T�����u�c�~B��X�SqB|��ɳzD�༖�H�J�D�(���}r��X�! ]T]ߋ&�������+�V `܍$���f������N'/�������t]�R�,)%$Ib���ӳ��/����:[E�����a �̓�s��|&	e�:>gIIGm�l��C!V"pT��q���Q%"6F�B�����`3��`t�CPj��s슠�d�a !4@h��� e����UL12!��V([��	̄��ĥV�i�+md���L��3��P��b���C���e�W�?u�E�2�DB@DP�f�-�f5���x��/b�: �s�l�ï����m4E+�d�B�ϳ�h�C �d�5��h~M�ӥ�<�ڎ��&,7�!9*�,)�B��>�dD�FUh�m1%h�&I����}�u!ɂ��N'9���1�b��Ȝ�\���!�J�9������y�u�� �(*����o�ۿ�[���G�ٟ��r������|:���o��K/�����������9K�����f�9 Q�`�!f�k����upx��� �o\����w�����ѓ��m%K�u6�/tU��z޴䶛c$"�2|�5X$�����;͎��R��!�u�(��Z�G�rʽܨ0	9�T��C*8����LOUUo�D� 9A86WU�f�Y�$M� �P���S�1� 4GUgq/6��>��!%M�P3.ᮦ?b����،��܏�����>��q���`��i 3Q��#��d�4����'* (��҈D@����b�X-�۳f6�@3siG����=�dH���MFu�,� �g��=x�@��>ƈ�nf%��S�����?i���p$0�l�!EK��l@��L RL�t���o���E}'����$��Di��(��6k����چ�(���Ϲ� �;n�H^�Ye�e�2ȇ��F����.R �����=�dɖ.e�Ai٭������ǀHH��s���ݪ[�>x�,�M��t�Qf""�b�  �33O'�m�>?;�����x�æm'ͤ��r�(��Z�q}dc3��~���
���0=�~�l�A	��>�e��h�q�ߗ˧�T�,܎��f���Y\ϟ�Wt�BԺ҈�D�HR�TI+T��TO�4�U5I�.����*c�,��IY�Z UȒU����-B�JHHL(�Y�'AUK1�d�`v��N�h�������������e�
byYn?���KV�,Q)�^]Q�V�V���>5FͮĮTSNV�T�FD�{�,�A+�U&ʣ�^�8�NB���l:S�흝��Qv��S��.�>���(�!�0��x�B"�)�&�H��_|�������?�����l:�,秧�;/��?�������g��}�/�7�LDT�r��"��$l8�� h׭�����ε��W^}���~���~px���3�N�f[��ۖ�f�k���]W��=����ef�9f����Q�_�Gв̖���XȲ��g�Kf;��(����YYٞ ��ziV�k�;�nn=X/�ݽ��7o4M#Q�	�W�E�u�:m'��D���#�pK@�ĩ�iRLGO����L&�wUj�=�Y�Fg��BR�Z�a�����-ǳ��cM%�A=U<S�H$#�MDT�i��!�V��CU�x��`�xħ�����lkk:���흝��3�s�"!*���r�
S��F�4<� E��_D�r�B�4���1A $�L&�������V���9em�ֻ�d���Y����䜬X>�sf���B圕PTS�*��{�x!�.��-�r�Xw�t�с�R��L[k{�2�r����n�^q�ʯ�ٻ#HF��^��`����Qŵ��D����eis�l�Iz�e�Nr��9���X��Z?$ND
��A%���ѣ�~�ݻ�ܽqx���X.����l�-�?���C���dK� �^n1�T�Z*�~�\ �o��o|��o��������h D�㍛7~�w�������?yrL�U����X+,�Ê�Uɗ���<ck<S2���PJ��xބOUE���F��>�O��FZh\�k+%��1��Jc}�SRc�X�:h(,��~hM���B�CZ�Ġ��ڦ�H�ۼ���oӒ�� ��]T5g%t�J�bB�U�~� A{no �&��IQ\h�DK�����EUE%���s�)�Yp��	�&A���Eǲ4����²H
Zs9D2�8�de+�6�*'�	u�֍���|o���,�
��"/������6{h����]������\�/5�����6!"����I��s��O�����>[���S�����W�W"����d2�Lr֔2j�Ih�.��5cF4��i��r�Z���~��_���~woo��������m��i�w]�]ۻ�BL1eo��)������e����F��EmJċ_����w��_����LIӓb
�Ͱ��� W�J��6�P���d&�u���� "��.����o�ۯ��Z�c���}??��}�6������C&�bo1ΜbJǧ'���د��Q������6���2�0�˩�R3���.�D�P ��R�rԊ�J0�|>�,f3Q��.ے0�HPh�&4�%t����ϵ��������������s���(��j�<\�9��R	�\����U��)����vww��Y�%怈N;j�""rpp��o~sk{���w�ݻc��SJ�2*�%�)4M��׾��o����'��H�=G;TUu��=��������}�b$"$VͪBM#���}���o޸����ާ�-�˼W�������! ��H�vF�6��j�h ֡B�7����b]yx����2�h�Xĵ���k6�Db"���շM
�������P�Ќ�乮��p.�g{\6x#5̢)%Qa���Ug^���noo�گ���l��������_~yrrom�v�wb�~iI7B7���1���窺Z�B�o|����?��-�����}�omm����dwg�����[,�?��|y�S"
M�,Ś��J� �0���d��P�b�H�w��7T��:�V����wj�cZ��hԑ��ڊ�`P�N�eE�Y���X����BA	5�=s����W��%@����r�OR;��ORò�����uGB�]@2�~�XUo�g&��ua�jm�8|�r H b}� �p��V�Z�"\$3��P%��������C�
��`[����hh=f�W�,��J6sb������PM�L)�LBH��0�%%�<qe���6��W�� '�$v�������T�9�!*�dE$f��K�������
1G��cv�:KF��4~���w>0�Ҫ4Dt�N$˿���տ�7�v�\^?D���=E�u�:8 0*��t�٢�O)��l6���s�fQ�1"�}Ҁ��J��u�5����ζ�>u�W�	$U� �nZ�0� �j�4aȡD�����t�f$ �7�Ɠ�
�X-�'�M1H��3�s�: �Ā`)���Ob�e=9���W_yEE>��>%&�}�Vq���{k�W�U�wݪ�~�������l���5��T�I�::z�R�)_�v��_�w�n��`�*�Ǫts�.���PE���R��y�U��� ���U1Yu���&&�qkk��3[.W��|�-��I�X �φ��H�9��[u�h�������\b����N��CU@3�r�Y���Ly[��\���@Ĥ�s�ښ���f��NT�J0P �d��)������_|�����>��D��1G��Qє����7�������~����}���#�O�`QUEP�ӿ��^�~=����'�ľ�L&���Hr^D�����ݿ��o����Ǐ��{��X@�XD+@,���*o�\�>\H�,Na��U�9*Gc�XUaSyc�aik�[�	0��$����G8p�K	���#S�"�*�����HdDo��n۶m��|�r��^D��������ͷ�\,��O>af� �ɰp��꧍W��t��$^�4���D�ӟ�t:������b!4O�����Dd�� ����l�4!%I)�ָ����f�U.��),T�� ����eR� �4�6�T-C�:@)8���������G�)(���t��'��3���#%Y��d"
d	�"��r!# d�}g�Y�L
��h/"8�;:aR!��1W�����YF/##���[�Y��)"Z���8�-k��6���B��3�0�C���g�9Z�M��b$_GD3ſ(Ы-�M�˥�9V�Š7���谎�%rvQ"��(b�� ���'���+{#Toq��2v���B�M�c��B�:YZ�	� �����R�Y�LkE͜sN��Hm�v ����*��Q�=�����ѓ���}����3x�i�r��r�q�Z�u�Ͽ��;==�O������ʯ��"loo�۪�\,����9�Y;⹮as��u��z�7ogՊ�FC�0WV��<8�@Y�}�O��EŘ���HD�0p B�/e@��a�X���6��@g5bɔ��*~��	���l�؆?��я~�CQ`b���}���<��ɧ��*��n�pk�u�}�>��]�q�f�N�����>[-WM�����WO�N�|��ɗ�W�,��d(x�����ʕt�
�5o/e��
�b�@�_AdU ��t:�LD��;�GDWe=���xVpO��ﺶi�& ��2!�9��iB�s�Tr�Y�E DU���,Ez�KD4몛/�sf6�R��3��@��ǟ������(*0s��	s�99;��O�?|ا�A�$�t~�B۶1���y�ɲ;lnM�fɐ���{{{M�������B���R�����DO��K���2�b(0��c1}lɦOٍ�����50��Q�\�g��We[א�%:`7u����o^����|�KFvN�%��&񈊇�������C�?�������}���}�����j�IM�!�֦8k�}|PU"���5�s��?��?��?��M�.�m�g�<����}$\.���ĔS�ä�5M#�L�}�1���]KP TS�P6Q�٣�D��=��$���oTUsN�����b�! �Z���/�Ḧ�=��U;,UR/��BW��P@��*�3Y��Y.���٢ێ�fY�7F�����[�.$4h��uQ0�3&b��	4O�6�И]���H
`�(mU2�f}�w��y]8��h��׉e��Ņ@�����Ge�Gf�j��z9�{q���H���G�7���A�� �  ��u��j%��6	�<i�� ǲ/�>vܭ�n�Z����rj~fx�����/ X��
j�7��W����D�J��N�-���6D�[�;���"1b���v:!b B%D���D}�M����_�%�M�O>� ��ko��W�r��=PH)=99��>E��6~=��*���U�Y������&�\G�B��b��aҋ��B�f52�hh����<��-"i\��J��E��8�����I���v�Ddo���^xg6�yew{k�	�s������?���ɓ��/��ҋ/3��>������wߝ�f�'��>��3J��dT_�x q�l�zu�n�+5@��_H�l"��J&�������)�]���\Ic��d0.�h!�Ue�\�������v2�LcL1�dY1�튙����S���|L� c��\���g��!�������ak{{�\��TTM��i }���w�~�iJi�u!�<��:Q4��|���?�s ��O��Ҟ���Ha2�i����?�я����7m�Z��R�Įv5��/ƶ��=Sc�8�ܯ2������)�����]}i�~��*V(��������� X����ߒ����0�;s��RJ�2�lQ۶�٬i��d�\���{|�a����m���ݜ��.�KS��s��Q-�iF]YW�W�|v~�b�L'&�b�V=�\.���B.���}h�0�.�*�����B;��z1O�dQV!p��v���v� g8��6-U��Ԍ��q��b���oK���+��G����P��h.�ҿ�Ĉ�R�Y ��3T��ՊH6䇭���%RJ(����#�eF�P��F���&�R'"#��*�݁1o���f�7�����Ћ�g< GT@TU� �����y����$CR�:�~Ԝ_A,�υG��$j�n������m�vb��17[��5m�sv���*褝Lg���������3���X�Up�z��7�}ӓ��}�Snڦi""�-J@%�k�{7���!PP��M��E��98CX� �LL��i���|�W^ٿv������Aa�\������J���߂�vH�.'��C�uk��2(�湄��V{���8��X�[m���P�ג���[����^#Y+�L��*�Y�`V>ǖ��>����&�f)�d��08�O�q�\��ε�sӄ٤=�?�ʯ���+���_;�v�p��*�}����_|�/>���G=z�o�t;4�g?������Ǐo޼�4�r��R��Du�� GpK=�cK.{>�UV	��~��6���-i�R;�jJ1�:����c��fB��q#9�_�Z����7M3��Z,1F��[�_ʗ9E.Ւo��o\J����Ac��d �dO� �ժ��� ہN]�B��g���ѣ�#栢��1���*k��s~�����H��^E�HUbVq��ԧ��ӓ��z1^t[ܜ�C��
a��$M�4�>g� Q�ܫfS������ס�# �6��)��X ���6}��e�:K�/�	^�� #�72b�����*H�K)k����:I9M'�o������ YV] ���z�9�8����g�=Ʉ����y؀��U��̈́8�����<����$��h�3�\�:Kޔ��
�oxcAD�q!]�&}K���w��.�We�}��ԄJ��k�j��U���U�Uh%U�,�j�G�������'ff��ڲ�ʒk�b��V���X�=D�b����%#$cE��82
!,�C��W k&� H̗of�TU�F�&�꼋H�)�����"���}����~G)����jX�e玞o�] j�ABA�F)���2�vĊ3�~��XE ь��-˶�q-�ɼ����AR�"¬ ��}�@�4�2�&��e>�眝-�-�z)��ö�l�%������r��ł��`/���3�L 3�����v8�;�ZD����2vۓ�l:�U-B����}Z��݀�Ə�ETr�:]�D��5����_~�e �16Mk��%�����lmm���/^Y"�i4���0-y�.A�?�&�~��_�`�����P����bV�mv��!&O�1�š��J�Ep�e�am��u�h�	�����!���>�Z�$")@�w�� �j�ܚM�g[Mh^����_���t~v����"O�<��޾}녔�w޹~�������~�ᝬ���_z��7�}�]#���2T^���
?����E��9~���Dfc�I��V�&��ɨzS��e���~������f)��ri��-e�B	����Rʧ����doo9�����ד�"���6�ZJ\Mr��dR�Ɉa�ʯ��;D0b
朲XW=�,b��M۬��6�jN)�_�~AU�U�Zo@�N&�s���qaC&f�����9�
�`Q���r{�P�H�@���g}#������8c1���@또���{�����}kd4t*[�]�����P��H���ڹDЁ�u�!]�9_78Њ� �����Tԝ�Ř����U"UsL��
'MVN���c߿��K���J�"
1%;�9g�t>?G���'Ƅ�%� �d1J�(>�(h�����e����8��(�7���GB�R��U`$ `bf��9%U�N?^ �5Ec�-�����a��͚&B���qp�j��Xk���Ʈ�I)c�B�o�_�JW��HR�))�kt$EmKk����u2�(@QUf?~1�1����Q�hP&�N�8���F�\��yx1FA�
���(��ޙ��T��X�]P+v���*�+&ׅe�r��M���`��z���S�l�K/Ī��f�Z�%y����Y#*�g�iJ��|N�[[[1v��*��k;&RI���c���tkkk�\���y�53�S!�V�b$�^@@�g�@�b`
Mf-�,���M9����O�����������)7�������籏̓&4]����$ �)}�嗪��Gmmm�����nܸqc2��m;�Ng�Y`���w � ���/�TU��O]cu+߄w�Qd7�0G~�������P ����� $+:�`m[oc/A=-M��%�2�ܵ*EC�ʃC���r9F��������͈��3[A�q3[�\��2!ͦ��|	�;����ruvr���Zt�}�ɗ_��?�߻v��'w�����'gg����W^�~�h���~��G��o��b>�������_��h��ȰĎ�\yY.f�K����)�Sf��!�fk{�m']���^F��z� mʽnQ5�(9�}� ��ۻ����J���T4�ll`́9�[A�'�l�b_X+'UrngP����M�a"Q��5��1!��!Ӓ�U%� ) �N<(�!XV��dH)�j1�]�l����K�
=U�9�!�R�^&O�qi��,Pnp%����"yeB&�R�1��R^�ZZ���EC��w(UO'U1/TUbL���
)%d��s5�]�������P蘐��d���j���X��O� L.ݷ�`�`��D��K75A�I��,��'���
=SN1F���.�䡿,�$�W�yp��ܛ��[n���]'��!ƘS��b����\�ܣ�����(z�x� ��p�
��a|g�u��8WSGTTT$c�=�l"��ö�_�xl��:U�>�i��`M9q2�n�n1( �Ok�����+���x!�0��i6��Z����q<]�Ԙ<\D�e��U��1�)�3DDB1�:g(�,�
+�
�HFQ, ?�1����u���L�xU/x��z�X�xm,V�N�/ܺ}�D���ggg���������և���L412�*v}�E��O9#aL �R�q#CP����ܶ��lf����/r�UT`Ff
!�M������ lH����f���?���w~���������%�I��]��?�y��/��7n���������b��;�RL�a2�"bL1�hF3��6!|~��{��c�7����Woݼ�����|��o~��:��������5G��b5�e5�W(K+�sa7,�BF�{<3O��x��V|���T���ٕ�󬢆�P���R.��:m�h����
�*Z�Y��FL��W`��6���&|z�n�f�X�>���=I)�f;��''���k��T����w������ݿ���Mï��ʪ�g�8��5��<]�����R<�]>�k��L�ߡ��y,�		�j�D��ɬ��if�) t�.Es5 ��2թ%JU���lH����j:�Nf�ɴ�1�hD�`�[^}Ɋ�?�hi�шTs��K\}L]0�H!p0������h��l�A�Fiv��Q�<�
,Ȯ�"V�n��ERRDjBB��/���ym��klY;�2�fK�9��7�
 PID��Y~ُ�����Ę<�� ��4�4��A8bn��%*a@#�R &���@��f��"Y��7����S�������W @	!p`f�Qh�a.M�lmm���}��ݣ�'�j����[u]�X,����n��Ռ��NF�E�㽨%���J$�~�0>;���<�!@����������Ǐ��12[q�V����V��4P����Z�D0K���+�U�mLV�N^�f�,��E(=���'���Z�=�2BKC�T�r~�A-�XKI	kG��y�>�c@�HR�kpaD�X+(U��z�	�Dƽ®qD
̄�@�G�%�X�y��S
!s2٢����eT[���SJ!��"�ݭ8��R�)�n��8š���Cq�E��>�;#32��֜��^���'xea�`�Z	��r�<)'�8��ɸw�]p�-�.F���:�,Q�Z�:��^�ӱ��_B���E����窮���y������z���Dwll�ۿ��uS�p�IN����!E��x(��?r&%�)j�9�c��RSӊ�YL)��>�ɶ�j�J�7pk?@�a����.�j��t4�)<�>�q�7���D�2�E�j��ڰ�g���S�:8;;�T��d��E�8�؈�k���(�ѹ=�a���y�����y�q��:��9��2a�PS�T�Ց�cW�:��8��h�8Үھ�n���!O�I$o�Z����VjVh��9E��������D�V5O	�w��i��
�^4�i۷���t��~�i���4*�z��럊�w{^�x�j5�{)&����X�Pr�	hw��"s�s���*Q`�����z=~+�~9).�s�v�||��|��?=��=��R�2@�Dv%���Ӈ����Ö��F7��#v;�k��e*@���\�����tXb��u0j���ې|d���}�|}78���N�D���DC�F���F85ߑ#�e�AZ�h"�>oX3�e'��M��E��2�����r�	F�6uN�-��7�翔񶫄�%b�� 0O�\��Z�����}�Xy��Z���	��0!�s���Q��<�Q�<��4[.K�7�npY5���<�U�[�p5���N���ג�B��:ޞz������ë���ggk�A�B�{]�?��y���=\=�0w����"ٮ���q26ٮ�|�I�<��ٱ�/�T/c��7><u��m�����Ǿ�w�-���Z���&�F��7����_W�n__�tVU�kwL����5[ �I&�ͪ;H�����`Zt��Rd��L�\4�p�Lv=�M.�O��S3��B8�W��d�.6��*��#���I \|��8��"�em�n�C%�sfk�Aq�O�Lz-�����dAe/5E0HI1����K7� ���҆{�rA�@q_^#Pl=/��mLz4G���\ec�g����k��<i�1��g��������
&Z���𨭌4jh�������q���b��	[�z����{����??/����T	-�|@�(�8���J��=�-.����_��k�ԟ�{�d��@V�(=�4f!'�)=~}���0�S��m�u+1H��̤Y��������ͦ�{�}W��+D&�2l	��)�C�V$�\];�\�+��]/n��]N���ڌ)�{���\a[&��¥;8mſ�:�7ر��tC\;K��<2���KD-�_��%hK�Ӆ�����lRDEl#�+������Q�p��ۙDt/ؓ|�ڤ����K�<,�d�ʏI�k��b֍grv�SS;::>�jl�8�߿z�	x�[�hO���35��f�m��h�R��UL�\Gb(6� Ͼ+'��~�9���3�ڃ��u,���񄏨�6=��m�QDt<� ���W�̸�/�l�Ĕ��4'q�oף��ul{���k��`��(~)Y/};S�cҮ���IP�S$d�5?>xw���7Bo''ZL���)h��Q<�j�5Oy�9i�>U��1V7���C�(���Jj�Á#���M�u���@�S_��s��	a �x�݂b�q]�6@����Cפ\�r��i�:����.��Ǟ�o�#�����j9� ����Ar��>����N��#~'P2��Y�:"�M~�d�K�V-��4ڷ�$��W� \\��,��X��e���k3�p{�w���uo��qSgY��cݝ��.������;�&L!c�E�P��R��h���t���t������Tsn����Ǐ������ն��"i���xjPͶ�(]��,j�i*��Io.���q�^r�N��%P��}���.�Pۺr�� ��ͭvBH=�hXyq ͹'�K(�f�N�1�#��;�E��P`�<���,(�4/��K�eT�Q�[��K��Bg�M�0甅
6�S�-�N�
3,tdІ&��D�(�hQ(��K�H�R�K��q7R�ֵ�@�RJfHP�U&��
0u�!�r1(ِ�rV��p�����uL��j�v�ȯ� �ޞ�SB�U8&9�~*D�ݼ������}ظ�*΋%T��T��������S�`(���B��e���g���� ��*W�����6��&�R@��Y8 @f:Vk.�,%���c-�1�O&˝5z�&���މW��n�`65�ޘ6����v��6o6szFҏ���@U�@�Q��׭,�qlѭPw;�x�z�1yH1x�;$�1���$��Ҙ%O%���ȀO���B�ˈ��ƨ�-7b�8��3E�����3�E�I�����M�(,�o�#��`!�yC�Y6P����h��\1�Uʿ��[F��|��֚"K���[gs���ɑ�Ñ�ɚO�'�[�x��:�L�Վ�29~~�v��)9'W�ֶ���*ߛh�����Abb�<�&M��wPpl�/VȚ?�M�)�w�Wa>�n�n(�w�UCL���vBY��:A䆠�˲�~ �f����ҝ�����F�_"cY^-�9a���'H�Z��A@]!a[��jW���������8����r�h�E� M�v�����P�@ZE1���<ۨ�9���;�C'�)�0� t�2���,U�pU���o�2�9���K[~D�4��oqk�{����/�do�+�6Ύ��ʞ�	��i�Q�cL�<����ώ�Y��"�Dʹ+�}6�!5��eU��Yv.��M����A�-6V�kZ���n�� 8n|��Pw�3~�{:$���q{z�g����4o�S� �C'����)���ރ&E; ��W6�7��>?11Q�t�t���U|5�d�����yq�x蝃��s��[+�����[��b�wӢzӑb�j���k�;S! �t��E?�!�������ũ*���!�n����MĄ���������é��0
���~ZM��Wsi*ܩ��G����CX�Ug60c�
G�_��0�U��*��_�e ��ǻ��s/0�2��b�"�5|X�w� �$�Z�`c�Fii�}X��E_#�KuEcra5���7�*Ό%a�ڬO�͔K���r��ڙ��[\WW���K=�N"��+���$K5aR{�^V9ƋUW��7n�\kv���|�8R[s�:`�a�,8WZ@����S���)�"
.�S�&CѬ%rE	�2��)KM �8�$=+Əe�$�lF{�`C~��	��([���$OQ(���~7��X�*�@O+��W�����*Q�W-�r���_���?l���qj��{��%��ɴ�b��GW8q�Rbrm��4U�&b�#2�j�Q�G��K("���k�{VH�������:o/�)}�#7��Z�2Gݻ����Rq7Y0��A0��VA>�u�#c��S�QC��O���bz��������=a�7�r�4�=-v]�͚9������)��(��+���T�Hrs��E�T����>L��,Tz�SN���w.�B�;WƌU���$�?�"c��{�Dۿ ���t1e�4 뭃o'sM]G�v��Wv�v̞M�,Y̯�JA��?�n��M�~��Y{V8ƺ�j�����Yъ8�ܶ�����Y:�z`�Ӭ�QI+=���B@�6X:A]j��K�k���"< .LX��%Z؂]p�(v*�C��Lmt�B&��v��D�S�qn�sf�#�gc��FFU�]`Ȣ���gݐ��������bv�(�?I~�)#�3�M�DK�Or���y��S���LO'���R��}���n �*r�i__[탫L����wA�����V?�og��'2�;�6����B­��;��&&��7�eP�[�'c;�RM�1����ß��8�ڥ-u9L��>���&LGs-O7:�z�HHs!�*�5F[�:�+M�!�Z%�D��148kj�q+�@��9�C�B��j��
X�Fi3X�\�%쁌�5݊|�p!�#/!&/}�<S�b�X�u��:ɮ~C�v]ڔ@��O�������?UDX���Ċ4d�W�'PT��?�sS�rщ_�%Eu؄E��;C�`r�"�����%��̋��v�%���ee7���<;͒��U��BH*���Y������А�8�q+������K�{�t��<Œ!�5kKE%�mゔ�hA��#_EK󊳓Em��t+�e)�����i9	��S���h%eH�4��?�f��H�-G��X�62B�[������V�'�/�f��n�u�6-)S��K��v=�zx��8������o��ڠ]r�n���������n>n��&_��W>GL�����Kjj Pڦ��c�`)U�L�>d�m��:�m-|},_�����+#�^S\�:NC��4��P?�������6m�U�ͮ���ꈞ�m�����7��?�o��ľ=V�~�f�S��u��TZ��&��HH{����&�mu�Q�ё�ȓ&��
�P���I�����	�Ƣ���:j�!�����t��a�kYL�ʊE�>C�?��YkFe?�撈�^U!!J\(P�C������(�1T��#ه�ߘX�2�8}���gkX]�β�q���´�D)�m*ܖ`�!��Fh��E~�nY�MtC�%���㥾��+������t�fZ�ȱ]�ڐEBU��,�X�W�W��jp�rP
`����*f�a`�L�O8>�͠����p��M��=���r�x��6��$��!�9	%>��lJ L���І�΋[>��Y!AA����������g6^����ruG�DͶWWu^w�>{)
11i͖��15~�7��]����$�����VP�E��nrκ>o_8E����t�0�'ů���U���ڨ�K�����a��~�?�髫�����dP��������aRI6+���uw��w�ռ�S����H*l�'^���%��_Zs�0��t�*:h�c�}ra�m��]e��@R�[����)4�^���t���_�8ľGF]$��e�A�n?)��}�,=���H\-��A��r+����Ճ��n�7}��B� �Q��T��!_00qM���;S��M����G֊H�����r20���wt��;k��eRu��ٙ�3�fy�^��k}�x��L�B�*z�ڒ��,�v*����lxW��<o_�ߧB*�Vp�c� �=c�ht5�ٞ	�de�B
:�4ʸ8x���3�C����+��2rb���2�@���P(����j��A{�5V���v�)ك$<��"z�9��4�)
_��䳉�W�O�=����'��Gd.9���z br���Y���ي~�+tE���PC?m�l܆���y�S��`�rT���f�eF���)n��&;嫔��1�_8���i	�S��_�˚�j8�b���Ȁ�j�{�I��ht)��?/n�H`��7���]ܩ��2�?^�k��G&�: `��b��!����Zi����j0�y�����|��mPḔzL�1ҘƵ�0��,W/�fA����]�8��N�HOO^O���d�j���_6[�"��컜�ξ��t�>U1�2V;9:\t��R���2:�T����S�咉���]�JMP#�Qu�VCP�S�� ���`m��Q�x��.F�؂S��9�w"��W`�� ���!���Ē�L)z�2�Kł��F��>Q�<i���b��`��Ts���������vb!�WCZ����?�Q
�����؟���:iG��-6�- 7�^�٤����U���}7e�����{�j��YjE�K�f�}�z?2{��a��0�e��4�mx���{^�v;{�G�*(((��������������#<<k�����S�O,�x��M]|i�?Y
m�L?��((���Tw�T�Cu�Y�T
����|su~}��J�誗�,M�B��o�xYб�xx�<�_�(�QDCZ\L-�0+?�1$�E� ���`�(F�7�@M!��7,yH涤����΍� /�Eƭ(@ Nm��K"� ���ĥɞ�ZJ�Z���jI� ��@ӕ/2\(�p��*K\�i{}��k���U0��Ct"�K�j%m�"�Z6���$�]���-���))dyj�AM�yŉ�Y�)���	|��LG]��os3x��	WWb��&,�$0��ti�1�Zqp���И��sڦIBJ�i�׶��'��<���,6fh�$�矔�S�o^#�&2�	1���'������|�������M]/|n��=�~����q�"���/���D�$İ[}��ì�(k����d�������+g��	3��w�v(��&�����8��~�%8���r�W6-�����Y3��2`3�%�dT4_K��rh� �]iĉ�F�ҥ�a�uQ:�կJ�{��!�M������"�U�����ۍS&v�ng�1���^����/��%R�L�fH���?(Q�vRZ��T�8�vj4��C�)�W�H���|��e�
m�hM����K)/�dV����&2|V��2��Ђ78���1D�g��|��.�n[
�Ao(��4N�O��5���'����mH;���H���������w�~�|��0�=/BV�ѵb�ˆ��(x��w��6p�d��tg<�w� o�WK��2�������h4Y
����}MVD��|����2��,T�	a�ɀ�"�~_�M��'F&��R��CZ��T�ҨE�!YGg�1K�-ˆȖs�],qi�K��{'�L4��-�Т����s������j4��5*�a5�q2@��<��B� ٰ��.%JP��Fjs�Q��fKY=���]���c㨅ݻ��4�����{4e�O����n<��K��^{VS�!����j��.QA(K�ؾ�a�}������N��Afք���5�����֠��E|�.�ﵧ���33<�V��zh�q�w�-y��q�.D�>�k����;�;������ ���$�i���� <����&�*K(S�-��d�g1�,xa�xT&7CP#����{��S����s(­R$]Ǝ���L�����%�שIV?��)�#5�N�T�۹��(	 �uUث�����>�p�R���%�s���,P$Ӟ�?��u��
̸���6��G��-�`�Z�f��o�d��cy9VZ���;���z[Rq��,ՉX����aFv%yVi��M�hq����H�����L��H�9���(���'�qɂ�!�����z�P��ª�� .8�W��XF�e���r:�wY�]P_��3�!;�eiG8 �������Z]{{Ƿ������F2��f��]�;�����Y�fc{�'���?���)'����Ɵ�D�|���14������enF՟9��y����~�qKLR��I=�6x"�Xos���9��Q*�
	��u��ٙ#{*��޾)K�=���GN���ÿ:��Ŷ+��&_E���E��!�&$�͉�b�����*w���8]K���UnЛ� PB�����(*/5�������MY����db\��I��M��;Ӑ�b�������JI�-ӡjw�XG��]�������l�������&aK������L������y��r�s�c�]�'����u����]��F�3=ra����}]�6�v>8Veې�����������_|��XA����|7���p*����\s�˷�/�i���@c��CH��q0cz2�Ύ1��u�o�S$T����:L)W#�ߺ�+�e�#�֞��&��K��8�g>#9ѡ��پ������r�p�y����
G4�~&ub��G����hM��T����IE�յp�����T�b8�(�)[���nǿ��)�%k)�?��롖�g+�U�Й��S��� �;=7G�VmYd�eu����F��I;]��qE��8�+G��Ɨ���A��ߙ��h��JTy���??�>���k����Vt�p�
�3��~$s���B�gn�p�"����3��&x�������՞#�W��w�vu��p�!��+C�s�~*��N-aHҦ)A��,�Ԓ��ʺ=Q3����0b0q�'g~{��Z���ʗ��M��|�?�ri)����4t,+7K#!E��[�G�E��2��@J���[�����Cg���:��=$ϯ�>�
����0����J-�6'5@��_D.���7�j�~B���E�j�m]U��28�����ύa�|�����t�jiZ��0pШ�d�H" d��n 
����W1��WbT��Sd�o�aXi�H �_a0q,� ����Y�3LY!�Fq�F>B\����\��@'�8�k���%���<��}q4|n�ON6_W��η�;τ���vww�68&��ٲ���9��G.��o}��6�w�|7[=�����T����X��������?H�jO��ݜ��͸�tL��G�|�[�=cPۣդ��4@J��.  ���;�;�&�E#�VNc����8�9��2����e���m�m����z-jw��f������(d���A��@�q:6�w`�f}ccÄM��Բ�L���>RRڲF������v��a7˾��c�����xzz*_��f3��_��FG� �����MU�H�15�W��Kp�S�d1�q;A��}E���m�5��E�B\�I�2)X"�7���n<���e�����Ҧ������;���vp���Ň�07�&=c�c'��0	1VQ�������Ƣ�w�{W���H��Q��G�����,.�1�bA�wau���|~~��,5$��:r2�/c��U�An�������=�tR�y�y�_��۫3[���7,&N?fT�Ҫ�8Df�/��U�u30�`D"e�u��"����fF*i��d,?4ao�SCE���̷y͔'hDg��>���<���CZ�?����7����outn�o��[qR���������1��M�׺޺鎊fi��2�[&6�ɁeG�Xa0�9�W��Œ��Ӣ|	<���K�8$�����noʰ���N�0��pŨ������tY���X�;�d������T����d��	u:�G'{�CXfR��Z*�|�Hcc+t���Oq��lm_�C!����ӻ ��~|ϋ�*�kjy������ƴ��yn�Y���On߽��>{��7�:��+���"��p[��uC�|��r���8D{Py�2�-�E��+���d8�̣�4<?-���
�N�g����r����
FĦN�$y�t�-ѩ8]o����Z��;8�yF"���������늫b�ҿ����n��
Q��Y/��T�<-U�o7ZQ1u�n�gN�5 �o>��W���)�)�y~>�����hi���0�q��@c\1��C�on�����'d��98A���]��?C0V�, �?f�S���vk��^?^(�4!�-	��<B�./�ԑ�G��}{��1�p��zۥ�)M`p�7���Bʫ$����X���O�ǫ�'�:Mӷ��؃%q�-E��67��G�D�:��廉J�Ű�{ʅ�]ܸZj�v�ZMS�p���d������]�ӄ��������d�|���*s1�F,��:���(K.�E�1"�N295#��;�9K��^,F5K��p����-	<�Ѹ�}�	����I�j��D���yP�@�'5��Q�n(U�����3��5�]�=`���_%J+$��_/��sp��a������d�{Ya�sͽ�ɀ�Z�uw��R�*��c��x���0�e��ڊ�zk��v/���z�r�\a��U�<ʿ��ޔ��X
������j���!�фC�V�ەJ>w���{J�!�.�䧍U�ܩ#���	[�t���t��������-����i��ctF]Ų[�Sƻ����z����5����P��z�ktZ��7E�:�{��q���{O_7FF̳}��Z;�x��o�|�N�b_�������V���zH�y�^�w�#WAy�
c��O�e�A�DR5����O		����:�\CH�&N���bn$f<v~nn 2DE��I�>5�ű`�"F�_��α�n_�
���{�w=����ϭ�諾�n���q���dO���m��
�
`��P
j-�77צ�F��5%�R�0�hM��1�X�q8�aﲍU&���x&�-p�{펵h��lQi�n%C>�lqb���3�-���A�������;��;>l��4f��ꬼ!0���]]��~+���-O����p1v�x���;VQD�Bٓ��+�,{߫E_������Ӧ�����߅h��׮�3���w0?�x��jol�C"���F�ܺu>.,66�E�RƯ5b)'���yy!�	�:���1w�v4�s��E�aP��/3�%�FWƊJܕh3���W�RRc �I�LJl�t���	-�c������ݔ�˼��z��O-!��5x9�|�~>lz�P�u|{M��n`ϐ���ы9�mٹe���'i������p=�����7��z��RE"�J"K����=E�
��?�=
�f�Um؊FBx��F���y�{�:}��H�ߖm�\3��0j�&Ǎ+��:�NŹ�����nG`�&s�3Vh�yϹ��������@ ����/+j)U��wK�k|F������G���4��^��\5��wر��4���x����
���,Hԛ�y�8���T�q�?	_);��7S���_�Y��
w��c{=�>S�O��C�~����%������R�5&� �|�*�n����0��(2������jU�CU���)`�C!��&�҃��H��$�e��L�a�>�	n&���~:�lV���^9y���[��/�8�Ohha&(^�"�yL�u�c���[C�m�˪9�	999i:m�%J3H�`F���+�k�zy|<:*�+�Ճ��:e��c�j[�7w�82=<d7�%�$q�����:cUg<
vP�l�2U_$�3j�-��X��C�LF4\��w7ޞ�);���P �-Z�/nb̈�o@STjЃ�2�!�mg�몏�e*��m4�khkk�����V�/k���۫e��O�� T��(
�ɩȗ7��O�:A
����=��WTT�+pf�"����?
�[�	���Zf���J�y!8�c��������/��knu �E�G�Z�KW�ԅ�b�Xa�Q�|�ݤ]��(yD��&g@�QE�h���ԁG
U���fs�*�`�Hd:f  �b�42D����W�~4;_dt�A���m�lb|�=�Ҟ�Dʖu���Wך��NCd����gԃ>M|���}�9f6hsX�M1=��LpPGe�,���z]q:�o�?o�!�����K��q�����!���6�4��'#M�"
PD>C9�7�3ZU��#ndw� �P��& ,Ds"#�� ��$*�	�P�l�}�����#���Y��ִ��ǔ�/�ApQ��^�ю`~���;���q3-ml��h�Ɔ�����/����IF&���}pT�V2���{��/vz�>4�)//G���ۣ=�y
6��ɴ�"��k[�3���tp�27���͌�uH6���8�����^2a�z����������p������n�F{2+Y:1ux��3�LP�����/y�4�`8�uPs�H�wN���iY|������##?~�x%�T{��tP��v����`�s�}�uo�))�a6�266�[���8=9���".��gde���y��Um���Y5@PU�[�oy��XZ~�}C�(� +�y���ʚ��TK�|������V0��Ї`�mꪖ���j/7��CE��P�&ꧻ1 #��є�o�N�]�^����&����"=��R �w���5c����-l�UV�~�RW�%�J-d�L�˰��AOE�B!����8��8�g��ApD��mP�O�gIa�V�*O�?�����,]�)�f����`'��R*�X�O���:W����)+�d�@j6��a=��B��+=��0��0��,J� Y�f��%A������0�9@l�wLd�)�Fo$�C��ORR{�4��+|7���n�����"f�V7��
ʣWX�4*@��7�&&&���R(&y��LY�f<Dh�p���R�N�gkNk��/,L�����*�����

��^���RR�0"0~"�`FQ����ߨn�U��!�6l\h\���54��i���f2F�1�������4�&�]ؿ=
2[�j2� ��
�b����q���ҊJ(�BI�3U���
�dHREr��vԋW�tt>����bfb�oq��"��g�4�$��P�%�3�I�����2[1W��F��_���֬��V��<�>�FFgI�1_����2T�"�\e�神pP	#X/L�
!��$�Kg/h*rgR@$>����jD�(Z@ f5T�����h��j����}�8���z������k~p0��W�U&�Ժl��-,�U�kSs����e�qy��c��i�`*+#+���i��9���������pL�J�!����4���HS,`��Ut�X��.����,V���|��9~A��E�(�(K���]�+���N�LC?|��kŵX��6M�( ʥ�b��sS�ЌB{N�K��lqbr��a�l6E?�c!�P� Nr��z�]���b�[�� 6��V�w��/�J][B��f�s#��|���.��1_��}�X���c��P��/k}]�X>t���MkAv�Ú�l:��0?�t0����8W���Y+���ʞ��9�ϫuzX��rOF�(�;㎝�.����(&3y&R�8:����y �����"�Qm��8yFd�ߎ�*BQ������Dqy���;M8��u_^e�����ܥ�����/x��WQ|N��=�}�9.���!��	/�MIiZ����=�g�;��d&�ߥ<�x�ˀ.���39�j���M�0��8#H%(�r1�4�S��䖩�a� ��-�t�=^���0��
W9	НL�~����0�7i�@H�^a����c���NF�x]�j�ۙ~��G"<���W,�-1�q����Guh�r�z��vl������|y4gf���d���m�UF	{�����X7�By{T�N<G���w��!U�YQ�0p3@��IJ��Mf}��+�r�1�$ިO�|�^f.�TO�*�z�4�b�@�~�����A�Kx*��Q�a�h�U'�d��aJYD��������L���� $�` �e��$�e��Yd2����	����* �Ȫ�͢�}�_	>��
�#�A�%��Y`���5�����I吪��ߗ�1ے*J&�7�}&ӐϦ�Y�#
�k�A&)aw|,����� 7բB@�XM}}}{sfs��n����RU�Eh�r�`lw��8��5�*Y���Q5AMm��Q�Ι��د_u7�v���B�)�4{����iE<TîQ����n�����$ɴD��C'w:�a�x��>��8���A�T4oS��������-Na������{4?A|Z2�ד--���$A�DT0r4�aA*e+�N?45�[(�9��
�����1���_j/�<LDG�SFAK��D����H�83�@΂ud�}�6*u��6,�l��KS�l��&�֖V&�1J��vJ���� h����)��eioo����Tf]�ߙ��go}~D��n���{�a1D�+nľG�z_K������M���&��?�}�Z��5�7v�S������jf�-3�si��<~rr0�mw����X�����I�N@��,���_]�%j�K}�u�n�#�/��#���l���|+⼑�a�放��'�O��Dy��0���+���خ����ʀ�N��%�,�W�14��C<+��T�����L����c�,��V��6w��"JGS�rwet||\�����d�j���;�hގZjƆ+��7�s�pjrrj||j�9|k�םr�sݮXkņ#%%%���@F&/�5�����k��P[u}���/�@2Mk���,!�Nfi�H��r��;Tg��5�^D�!<�9E�Gטо���9?$���O][_:^�7<��"�6'x�qq�bHZ��|����<.�9	cu*nͅ�N��t�}�tVu�҃���zY,�V���MB�"�"_���x�qy\=��͛6��#$�JjÐ���3̾-|�џ���jz�i��ι.ta�c��U����(j`&��6m���00�%v)�2yj��o��a���h�v�U�2��;�m�z�ȍ�<��N�+�D9p��*&9)���U2g��vI(3_��vx������D�%�gr��ھ�Ҙ4�[v�F���m`X+g_zaL@ពī~�~Bݬ�@���,h埃��)I��,Յ�@n$�V�"�B�ҩ&P���b}D���̨D�� |���d�E��=��<6xf��*��L�]��
.��F"D�0���"_��[U	��P�՛odeI1�pW߼i(��N<�a��d��ϳ��4G���j�kg͓��l���
��l�C���v���La]���S�/��(���!>�[��%���z��C����q��7�Hg���]c�V��+(M'�-����~y�Σ����矂q� ���$r ��]΅+��{��V,G��HaBY����eҢS�:���d�&�޲�d������*?bϿ��k'���Y�������������՛�����3p��� �:���?���u�D,RYJ��6��`.ۡZ�xKh�B
b��D��J�b
�Ì�)�`ЈDhR�O��+NļAHOG�FT#��1R%l������ߢ",fǂ��];��(у�S/��oБ����~�5,�ٸ��@��k~��x��|��]����l��	SC�X�d�Nq�;s�,h����q�}X�s�!M��N�Gv貆���o��I�����>���y��A�f����r�<P������-]J�z����\��I����?�%ҟ� ZE��U�SI�Ѵ6�̲:֢����00�R�I�cDR��/٩'��3�/T�A�41v"�������y*5}ۉ�q F�������uH��J��L&HdQInH�Pʟv^в673���	��>1c��h-X5���N�zz���I��,ȉIj��r�eyy����*VB-c3WWK�"�3��"��y�(	y`��U��B9�(���OC��� ��y�D`��r v/g���c>J���f�����F�W��֟�چ��g�_xm|Yv�ֶ�7GX��|^
�>;���߭ͽ�̋���؉cc�p��q/.�q�dؘV�S%#ڽ�&�%\N_���`ŕ�Lǌ�a�z���L�:%��s+�C?�����ʦ��UI��}��"��"1/����Z��]x�P,ɝ)0�;sj��H�uM���0?7{�'y<s����Dl�f��B�˻(�Th*E��+�3#�ARM�̌�Z��> �X'�؃��0��K~j�4�\fCr��y<=�0�'kq	D��nH�h�i)샑����R�Mw+'�|���g�uq6I�	�ϐ&�"��޽���(¼�P�4}�v�B9ryfc��O��\"BSn��1��L���V��	�>�M��X����¶2wLLPJ�
Ϙ6�U����o�^�B�ˤ���)<װ����́�@ĝ��a�: ��3<,<���:��[�\p�nN�3�W#��$*�52i�ˠ��J���e^���֝PΏ0�~�,��{����F��8�������2��U�gn��U[
�o��ֻK�X����/��G��2,(;�څ��g�^O�L�dN��w���4���n� �k�h���oQ�˅rDxGI�|ܦ|,r�i�`�T7��q�"f�xbF�*P-t���Cə/�a"ɛ�ݠ.�^�l�+A�V��Y4������������Y��S�s�Y��+R�a:aEr�Ȉ�ÀB�L�(邺�ר��ǁ�űѴƇ�,g:B �a�,ݾ��Ih��F.M$�|�^l/��e�W��\���!aeDdxdQ�	���V����u�=�Z�]��bH������o��x�LN7�ި�^��H��"S�H<fҜͭ�ܼ��^�y#Q�^ne���wd�N��&įJ���o��ʫ�����h-���<9�)�{�c����s�)b()�Wu���`���aN;I~oH��^�rc�|��A�;I;R?����G Ht� I���c�8<tVe��/)Y���*]p��0V?0�<��������H@
X�J~�
�e�a"g��d��֢��k�Ef�"��D7�sF<�w�iho�������h�|z�*� ��%33GYW�GgeӅ�EQRZ@@�;�nXJ�;�����C��s��IiXJ��ai�}����y�kf�}~�Ιyf�&ۀJ)�u��4xH"�t<$���Gde���%z�9��BᏚS��0�
��:�,�o�&�9��Y�Ef9�Ӈ�񭊹l(Vb��:7>'���T7�r݌/�P�]\�ThX#Գ=��i�"��)��U��I����$�Dy*!��:�*{�[�a����$���A�d�Eu�T?d|���9��}���u���h@���W����g�KAa�Uν0����k� y[�>*��[w*�[C=�C��M���̣$r5�,����\6S�����[�?=����#���
*������P?�wO/�f�j1�ɚ��Q �����ER��Lk�Jv�i<�+���T���|��\`
�\�GmP`�U+�_�"j�N]��G��n��h����}$g	�}Ƃ�̛���;��?�t��A��#S�1��Sji9eS����#:3ƅ&0�_p7Ρi��ۻ�!K6Jd	��ʘ������$��S5x��Z��B��QȔI���Qȇ�󯂛����ٸ�h")�>����{��vn�G�.�(@����&��mݬ7/2@�`:?^/�d�rM�g	���pf���U�X���n[�t���|�f�����dt�Ӳ|�B�(0ٔ��/O�W�7�[J�����!��`�_֦�bȩ�͒�8�d��C��wg� ���M����u��:��mV9�ϊ=į+��yɡ9kb�%��3Jbe�^�,6&U����8p'a�hf�J�3y��{��D@��3�K6��3fg��&h�� )NT��������ӽI�L��^<6~�,����k@Ȓ�����5�%o�h��da>b767����$F$Ή���WyDy�Fw\9,�*���ӎ_d�U�YnV�Z�xZ��&�[i͕�R���Z?˨v��W�)V
D���ش�
��\6�y�'���9���R�0
�J�%������-y��]�l��M�
�^�y���<�������:4�����\S.�u�� �z9'�j�O��wc�]�Z��b��)S�ʥUQ�-C�)�KNϩ�7�$y�t-GQ4?&3	���p�%����֣����-{��V'����n��W�]u�^4.��y�JS�	���Ì���$V}��Kԡ�U���^[�
��ж���T�}�]8=���On��:���?�<g��j@M��.e��%��@�,WV$�	N_�Lhg_��dR���C�<Hs0+�,	bc�ޞ������N����ȑi����W��ċ�l�&�<Ѡ�����s|���Q˂P(רg]��u����N���o
Yl���|Ąyx��$=���8i�ֺ��,����2�� ��Q�������5�灄˦��z�F�7�!r5Բ\HH�|V���테��t�?Y�1�x��� ��p6�Cm8��ײ�t/�=�Ph��ha��p�SY���R���(�ʬ���_�K�}U����X]��^��P�#�������IℯdZtN�z1x�ئ����B��:��� 26�r�(��l"'��=K!^5p��3�1"
`Ҹ��~�w}��d"�63����z��Ԃ��V[ek��1~�ĸ���g�F���{����}��JҎT�^��2s�p�!5J������2�[GGQ��.LdS�z�1EpZifOvC	4��n A-�{�������Y�
䪁l2)�[U'�v ST�ӥ�C��Q}�6j���LI-�Vʡ��X�)a?'#������bQ��/Q�^
d�y�,Z|}X��[�yC-�n|���Ϟ��Б�Y����/�C��lln�7�Z^����!$�}�ٴL }�K��#�����<�׳nQ���xYZ:�z�KX6���Q��/�Uِ_�ۿ��F�[Y[{$�Sjru�%u��x_�*I�	nHG"�ct�"*�o�k���a"��ŏ��a�>7�Dei�rj8��nD���t��swr�Pc���rx�f�{�����=?�c�AbZ�~S�k��彉6ޠ��3���wB���߅��ua����AU�+6��y����:���������OJ���%�c�f
d�R�D8d�����)YX� V-��cᎏ���{�yl�z� �~kk�tඛ"�\����h�ϥUҞ\<���ɪp��p���~��\|&o�Zw��n�2⋿���z}���
�>�,��d@>��>u�ۚ.�G�U�rNy\�6O0��V4�@y;Y���(6��x���\)�;'�:�*�/q�Q��h�U(��`�6�G>�^�:��jD �*��/�C�W:5'�BC1�A�>E:���Gc�d��l�=m�f�t�RTS�8P#�ы�vjYq�3 [U-��O���dx�Us|�;��.Wy�-�$q��%�5~D�e�BQN%i穂)�J�(����� Q3ì�C(s���|{x�BI�Y�x�¤H�T SN���ŕ҄aȲk���#�ÏzѮ�pwoxې����4N�ϓ�c4�����đ"��������W������ i��f�t�Qn�h3D?����~�=�_{�&�dע�־I9�����TZy!"���A�A��CM.��[�̏Շ�R��q��y8{�
�?�kZ}���r��z�0�}mi訫�>��,��ݽ�B�y���mȯQ^S�C��ب�/b@�cJu1�o�^	�z��TK���4�d����l���-�4i���xW������Z}�$O�8Z���]!�8�<�ȑ����a�5E� ��O���X�3q��ſ*�꾩h��[�
�K�b��6cm�Үs��Vr�l�N}O���f�J���#��H�l�3��U%���8�J͡��G U��D�t�ԇ���ޡ�]��,�ʷзu50S�g$	��JLqG �d�Zn.]Q��=�^���g-sL�LrM %�Pz�1�K_�W�V��Y���U9u�燸{Ap��u���ji
�M��f��c�P���_N��G��x�����0w㈮�,���qlm-�)��O���
���ܺ.���̡����\�����+���%�	���<//� �8��ΧIp��c�-��@e*�=d�شRɖ^z�I#��{Q��y�������G��F2]���4�Y i���[	Z�`�\�� ������%�a|�.h�Z�ӡN��W�O�^��m��Ҭ8�3F�H�Wb
x��1R�Nw��Y��r�WK�3Q���(��>�v��#�:��p�3��.��a����w�"5��'(�t��k9b��1�$��3�����l��c�
c$	�5"?2���it�=+`��fHE304th2ps��Un��韩o:��F���g{+ȃ���(�ߋ�%��z*��>Ӻ���l ;�P��˵����{�f�43�f˖[��H:G����ap�u����@]�g�5R�my��M]{Ye���z�V��q��y�A�؟�ow7�\�Ѭ~�kG���Π�bԒ�<���31hmI$�z���� ���-h[o~����`gÒ�X�(--�}���29y� OOO��O�H�d[���!����q�j��S��� ���&)�XXYч����
��������]kVͱw�L8C�=a�4�˰����ɴU����uҸ'��ǻ��������/�����`�I�*����,VE�}y�z�I*����I�Wt4��K+S�G���.hf����Q��("�QL&��8��|t��K˫�o)gT�*��Ռ�)$�v�,..��'#������`z���Ӑɛ��j�xLʑ��n�Ä��1j���$���n�� @����!.\��2y�G��!QT,����i�0yb�8*E={�6��!���!����1ر���8�=&�@�}�i�
�xrQ!ᆮ.�S��u���\]{Q��,8�=)�hh�Ī���	J��eA��������c��߉)Þ�5?�X�ݱ�)�/w��'���,��:ĚSGT�O��PS�Oq:�J=j��h@U�v�ؠ�gn�.����	�j����/�J>�H���Qk���J�6#��-�(��|8Ly�'XiG�u���#s��"�D��#,b�⊢�y~U���Be��c�%6zC�l����)��>l���^j��k_�#��̩+g�fRH�V�����	|ץ	:ď��1X?\T #��*�Nw�����<�FA�WKXm.���ô;��B�@?���	do�K��6��<�h`��"�ǉB��OP�B�U'��X�us���wt|���Ai�KL)W�ɗ!8;�m"ŕ֫0�$۱���!；'�6820X[�	F�ys�sD/�R$d�xzj��Z��d��rf��1�23?��Y�맷j��8:9���PϜ�gi]����⫈�UX5|�-�K���{�g�?I��,��@\�dt]el$��:�C;����,�m��x�&Rʔ)�:W�\���h��>zXy�� �����5�M��)�,��i[��7~�R��n&Y�m�R;&~z/��+5���<LcVx��!ɬ�=�=
�<Sɀ�`lם]�q��G���E�Xi�s�!��%�|K�zY��k�^���Vɬ���Qς]S����m�����#�;�O�ĸ�i2��0�A9���2n��ZDU#����j���?3|��B�3�C��|���Sd�u.8�������';/� ����J)ZVj����&�:T�X	��(��-%�OV�`��;����<�o�*<��Ë���	�LML�u	��]�#�PO՗���`ͬ!$�r�c�|�' {��.?�i�^r��Nf�IkSWn�����r�Ȓ6��L����S}xu���v�����}�"�a�˿�$�!Ѯ�5?_�6�m��_���U���������@$�q�WN2��>}E�*��X���(��D���2,���18�pB=w�(�]5.���5z�$7p$����"&MFɴԆ?,�YGͼ��,�<��:�Fnnn<��Vx�3x��֔��`q�FEm����?W�:0�e�������i:}��hA��eM��T�:n3����RQn�Ù�0>9�G7v�?q�
<��çb�����Ȕ�����H�*�w��R��*���\�l��L�7H�$��u-��ߢd��uAVԻzlX��vxUq�7991��I#l�E�y��j=R�^��ׯ��£Ҫ��dǤ뷲Y%,,,5�a�i*d����	|--N�]MMJ6�j��r��y�zz%n�89�p�Zޓ���&U@��P��+�a��j]N�$gO�)�o�X%���&*���Ox���A>HA�<�S5���r�	�DV���۟FZ�K|�;E=Ҽ�ym�<� ��P��f8ګبP��Q��8���M��}�<N0�~��2A	�o�xHj�W�5<q�F(?`Ć�'ih�F����)������J���K4����;�Ї�rԨ��i����?¦Nf�����:��W����x[�/q�U�8*�s�I�|�A�ܹI_&ϸ�y��h����r=f%7y��6�Ta�i*�~�F��n��+�s��Pe��L�R��"�-@�<AGG�Y���e�_!�\�s\�>\��6)����gx֧;S�0N�7������X�HII����(z����Ѿڜ����ا���`wC]�k���$;Ɵ��ic��0��9�9�����Pf����
��k�O�@�TN^���`��6ʦ�s+�(�x��f��CtΒ��Z�l3� :5�mRo����8��cg[��	���II~U��Sx!T|U�Y(��߾�����1�2,h��������seL9e�d��q�g/W:�V]z ��>������"X�_Q�"�Z�]<���Q����S�����#���hr"�B�ƞ�\ 9J&�9!��N���r�]�({C,t���r��OC����׾��W�V�ST�Q�j�Z} �ܢ������Yh�^��^0b������+ȏ�x���*Ex����_�aϋ�C6@���奥;�<��?�g��k�d��\<<=--�	��b������ƺ"n7d�l�5��n�۳��m��#=>N��Ƥ���NZJű����"����2�NxX�җ�9!׋�9�t=�,={��Cߠk$j��\�O��2m�i�sݾףmn{8�$�V�����7��7.��<l?�ު��zqk�@+�q��+-�'V�@����̠�����e+�/;N����mm� Щ&+���a�Y�{�90ώ{���������U&�[�ۄl �[�XoީE�h:۹k���y�}�i ��	f�yXL��m�^�����X�h��c��x�d�2~�  @GWD�
K�� খx��g��&�9!3	�Kx>Kȼ+!2^��,��2F�е���,��mnܛd��[�ry��Y����lԟ��k���iE��)����p���FE`��� #����Iq��D=U�i��ȹ��le�_$?91�������[��gp��<� 9���a��y�{l��'%��������c�Gs1�M���0�ai{G��&%�z������ȣ���Rم�\��L������	��Ë��t��H�0��"�J���j� �I@w��7 E��ua�W�����Lq�~�2E��r�(r>�Z��:�n��ۉ� RwQ�@C�^��ۆk5�^�hC������Ss����zW��/]�T��-��Hl
�ᢙ��f�H�[5F]�������֓�=8R�Op��&Yd�3����m�"$ �e$�����~�0��|�gZ��d��%��EŀAK�jZ��Ҧ* Ϊ�s���i�A�%�)�Q3�mFR������Ap�d��
���)P�]����k���T�[5�@{�)�/�mo��ģ����[@8N�z�nW�EI�"�p-��zMM]���E��J!�6��Ҫ�,�)�ASuf���+���{�*���bb5�dr�����U����>�"�M������dD��y>�V�c��_s��D�S��^�^nn�+-���I?��������ɴ�TҖj�hT�� ��,���ԥk^�����'�ꝕH����x�)i����s��p0��GH+���T����hB8�z�WUnH�*���R��z�~夅������Y��p�Z��&�Λ_��Gq�D@��8��6
j�:�jG���͏�^4�x�.�X���_���mp�#�{x[�j�r�VϚ��n��&�����Q[!n�����FҠ6r��c�G��7d�I��l��+9GIB��u �.d��X�c�L�K��w�btur���*%�@���AH��fD\\����b��4���N�h%���G�Nw|�͵Qbzk�>�IhN�~�ˏ���u�������g[���Q����i�,<:�Թz����]�CX.�� ��/����k�a][]���zt��{�٣ss�,��H��l-hV���e1�`�\��q�#雹䙴
X��:�����)�����׽/��ƈ8����~�+B6����{%q�n�Ӻ�QF����;�(����yܺ��C�Z��B� �'�,���N?���6�<b���*ǅxxx&�$�ܾ�(W��Z+���F�#$��=]�y�=�/c��b�f���-�=�x��Z���ʑ�g��Z�4�M��[�m�dX.-5X㺺hH��?�,/��2�k������<���޷P��;���+D��i��g�kp:�`]댨���
��K�,���k�]������d%^��ji}
~n���i$�� Y��%��*)��i��5n@���?^õ�.�<�.�U0�6�2�Xuԫ����p@j�j,@uKv�Á�W����������!�����O��>����c�;��f7���������ߊ[��MMq����[��!(�233s�NE���ֵ`��
~��]�X��Œ �n񜃘������
|�e��d�9�9���m��
�r<���+&Qܶ������Tr���\Ѡ�����]HX��H��%kb
��|���{
r3}VM���	H�������6i�ۀ�$!ۅsYw�:A��/7���b��NON��\�<����qq����Z�B�l��o��~�TV�dJq�:*/l}v㱓�ltUҬ�_�l����\��/��]�Q#�Sy+���4������bM���6��/���P����rN�����l���Y1��A�_��e�'��"侧o�F	|����#E}}~����͜K�[����o˭�<!,���R�L��s���$Y���=��%N'�$��*��-F�,"xC,�,�Gs<+�[>�*���0Y�ԅ7J��I������G������#�7�x���%U�����l{R���5��v"�^O�`�a�F�?T�ꄶ)��~iv68�"�c��م;�0
$�ߨ��e�m��dg�/Ӻ�IR��Ŕf�DwޟŐ�����(!��d��T�Lc�+l�7Ⱥsg�ট�9��Q��,c_H:��[]D[��,��M�X1к���!��h_�xڗ�<��r���F�ޗ/���,z��P �b������& @ps �b�*A�\��I�L�(=<�5\YY^�u�<��\�aS|�.�v�i{Y/��=��N���?��9>����Q�4n��heB�n��&0Щ�!��M ��@���\2!m�6]V$��a�r��ǡ���ߺ/�����}�<��p�͝n�RZ0Y�̸�շ1���{5H����\q�������t����f�ͮXY+�w''������q`䀩���:��,�1ة�v��ӄ�L%�*x���ZًOh�3G�HM��*\��fN�%W�;����v��\xUW�'1o�'��O|�_)Pu5+�~ཆJ���W ��gz���E��*�gr\5R$�zӡ�1���@vVo�����`b�����eV�N��?������?��N����)#�~/	*��%�����l���ߚJ �o�/�BC�wR �I����o��Y���L�H,G�r�HX�t_�q"'��ƄD�B��k�"X�ʡ'�8f+������}��/^SA}��y�@>S��,�����<�%��0�T��_���LDq�]�����"������Z"xI�j��G	
h�v�n# �L��C=q+��B�˦fݯ�f����E]K���?x���r!�-C5�6�^Z�����:H$z5���h�\מ��H%_�c�HGt'�'+�h���z���B�.� AZ<��D��aN�?Y�ȉ�6���Խ��F��{{{���_{C���+6�]�Y�q�ɥq�,��E�9�ɴc���t*��S/�|=�<��Sza]��D���*��Trn������i�p�f-|��N��y�p��C�dJ�2�.9�?��4եB���J�M�����:N&  �ɑ����r�:��/�>`�1�Տ�\R	8������ �L4��]�E&��I���R�J��S�1"D��`!M�L��փ������R]#��F8H�ћX*Y����Ů��\N���/�\��#�n�,Ju�D .��W��B�贀9� T"	X'�H�v"�����n�s�bM��{hy)`��Hwo�7i��q+�a�x�ԩ��e�*��uuZ�nƽ��{�@E҉o��(n7X�m���K�+�]���g��[��f�<�������� @�L%MK�k]�Jmx�*��~Sd
e@�a���.U2��/,c��~��9�p2=;�::4~н:>9I��4��B���6"���\(��G�6%�H���b�{{�����f&���-N������/���[����+|��<;�G����nVNOa��.
�"`�`Z�
Q+u�!�^���ί��=��m&!(�1��ĥ���=)@o!�ܛ���/�Fx����o�ږ�,��sQ�T�Ca��]�^��NVV�g�!M�X(`崍�ON⫛�]"�y�^��ݼ�nq�+��hR�����{�"�	����ݑh1O~�M����Iw���:_[?~w���R�eK�ǢP�fj�~gw2�H}!5�]�����E�b>XM��VaƆϯ�� ����R�R��UcP��z|(�<Ŭ�쨤2F�t��KEƖ�����R�7x�k�Z�o� ?���报����5�[�p?f�i�7M����D	PV�!�T�o���/�1��H�����"��>%W�����v˼S�G)�d�/D��=��q�ݵ33�j������4��u�#�ڧj��\=�r�JB�]�}C��Axc�e���OH��
���31�k��"�q����7.(x���of/'Jaj�[�pZ�܏XoY����h������3�4����޾��Md>PZ;��}�A�+2k�5��;8>!��  P��
✨]_��w����Գڷ���'�2E�����NUTƤ��	�\�b�����?��g���2-�xx��h�U:�������O��:Z*���"*ta
e��;�W��������]�ī߂���=��9�L��m00,0����^����X�Ck5*k55��5�boN��+b�9�,Q5��:��ճ~+2�v��{Z��Ƚ��:H��<��T��撷�}GeC� ���9���������{_0�����wr�	�\�z#�&����v~��j��sy��մO�����i9n{8�����c�3-��������Sly	1_��9�:�Ij��ǎS�C�'rMI��Ϡ���j����E`�V�� ��)Ђ����.=���`�=�65C
�'����^8&���'j9:�l����du�E�⪵��qM�W��z�^n��h�n��=�8�x�����|-5E.����Z�3|��ͻ�r$���1V�Q6�#���&,�Q�ǈ�.^ߓ�b�0P�f]�v�ړ{�mJG��_�>������5O;vܘ���I���`U+���� G���;::	�#WY���bn�\�N�$a�S2q�c��'ÖA��kFzz�)ՓK�?��Kᥥ��?i/�"T��ŷzi�-����f��
z����\B��VW��n����W���Y����Bq�nO�p�x����²��B �m�n�<A�KeS_D�m͎ÿ��	?��c�H�̲�d4]7���|s�E�����e�_���/�j�\% �-���(������~*� \���d��Y=��|ꏑ)���3O�l)�]G�YG�*�����ܑ�gd�f���	�t�����c�m�
�t��Q����t8����x���i����x{5���P�d71�0�E�.#Tdx]8:R�B�n,p�ؑ����9�����T�gn��n/���㆗���y���v��{i*m�"b5��ً�wS�j���nK���b�� 5}��a�����-W�^�|?8d��o7K�uo�D�Rm��ޫ9���j�{ÀN��lc����H�n�A��K( �:�dF�4Vç-n��P"52�v�s�+��l^,�aW��s�/�ZŅ���:��$ ~}��B,|^b�S��/�3�Z�?"�og�m,�����zӍ�<�)X�ktc�L����5
�w��_��Ņ�!� u���O*z��>@2�8�� ��)��6��;|�U�-: ��g�ڴ4!�[��]�Z�4?�]4��M�\����sh^���%���S2�E��̮����E��l�������{�~9�_�.s�3l�ů�n㥳NLN�mB�!k^c���q���4�/җپ�r�Tg�ƭ$� ������<�/�
�Yˡ�zv�_��o�<�xu�2s?��K����v5Z(�$M̍d_M+;��K�{)�*�x8���D,���#�κ���91*d�\H��ove��A���es�*7�+<''����6���)Q���p�����ê�b�!�4!�{
��f��0���$J}4I��* �\-l�Z��k��h���TT}]�q�U�P���rH���K.};7ѸU��[���j_�$k���P#��ɫj�c��&t�xxI�����>�eg�8����}�C������_��;�'���K���UD�7"�}�&�����t���?om���iO=����SG��#��f� ɇӁ����=�'�H�N������9��ty��_�U�i�;����=�Ǘf���nzb�ߙL��#�n�x� �s�48���l��K5��&+��]����;����ey���8YsGG��D�oW{p��8�)�y�Xq��y'2� ��)X��3���1�eݶ1+���/��� n7��t}�h;�m*�d&���y-+3�Xߐ�\����K���׉���<{S�O��iaN^:��z���o ����$�	~Y�ee����NDĝUCji\!�N����1#wmG��Ԥ�~�i�x:���){%��5���J?���.��<�� '�_�G����uW�ГcXܥ���]����eȡ�{@ńrIt�{b�E^EZP�:4�.Y	|�="���J�C͍2�gH66�� �o�l��p�qvq������3@���r;�jsE��7����M�iq�~�@U&l�;Wm�]FX�.j�J�%'��$n�*w���(������K��*�%�`�����"�[N�p��.P�<���|����:���م�T�޼�P=�6{����k��J�B��q NR!��'��f(����qʯ�A�ƽ�yo��Iu`�'�4�� �|�jR�y�^�te�і�a,�������`n��9�N�c��<��S��lb�Y�+ű|�о�K��#��9��E9k���������FΧ70.>�#��y��ϙ>O�?׏��lw���f��a�Q�R�/N�
�>�M�yX�q}zeˤ
z~�������6�p��vkhPe�x;��ivlY�y�I�����rE|.n�����r����|j��k�9n�H���Rk�?��5���K%��ZWgqZ�Fl%�����E�ai��
�C�\q�n\���e+_��ϺWW��EFף��>ۑ����T��^�g.-�O�܎���Z�J�j?Qt�^Y��]"d���l,��谵�����>	QR�Q�n;�E�0bЭc�XUy\�s�UG��ր���1#'1���A��w>~��?��%���ц�tѺ'�{���l��zx�w�C��$��1l�vn�k����p^���1=�^	i}�|��8�Z��S��_Nh�l��H�G������#ۚϕ��f~������i��p�K�P��ɭ�˳r;>e����}\��F�{ēBb��g�!
z�jsۓ��Y���//Gs]A�~�>W�3��=>��D��Φ��N�\.M8�Z�L� �Z��7
�5�'&23oxT���.v���PS�Fg���1�/R9^.�����z.�4�T6c���=]��h�}���Yc��vۻ��y�([a��I��X��?��y>̔(�;Cɰ���~���v��lz6~�v���� �D�Ň�SWw>���������~����������l�������N^�nL� �R�r�'�w����|q���5��+������/B�����y
���U:6[������׫k��L�*��?��%������i�gs��	���UtH�gS��,/-q:�t�I���	����^
0 ��{ Y���z�	����Ѐ��*�Cbcg��Q��<	
$J�����pl����v�`
��j�]�z�g�P�K�_������P�gK3"=XSPf'#�c�s)�X�3�R�3vM$`z�k��.��L4�(�pV����X�m�|��ި�����SLcx��!2�^^���>.rQ�`!�z����%Z��'���˾!iİ�3�H�q9R��L�a�N�r��Bk��$��Q��������wPj�[��'_���Sc�h7Xzr�1�&7Eh�)�/*��wKC��RӶF �=��3�32r��v�f=�ہ%<;>鷇�ƅr��U���u�|�hИڦ:I��&�z*��-��_�|\3MQ!zY0��cyi��Z�b6.M�9��4��sb��S��پ�(�'��i�NЇF�]nPZ��F$G�h(�'`.� *�H�;o��]���.��}#���G�C�
�sR�'�%r�poD�a�+JD���nfȳ��Q%��+�/�?{�moꥏ��a���[�6���6h�F����S����YVK�P(y��O�q����u�uwg����A��9������"8����?�������͊x��
vp_?���*��S/��M�V�B{�Re�|{�����
΋j��~,��&Wܸ��1إ#�3{����������Ȏ�;��̈@Wf���~A%WdɁ�˳9q�3�!�<(�vp�0�E�Q㦀q�;ǭk�a�z�i��81~����dY��Y�ϲ[��`�MMMs����nkN|�;��]�b����t1�?��Nxs��k�֜�"�AA2:�xH�-�1|�7���&R�̗��NgH?���Q��"D�Qq<���F���
��I���u�ciM����P[�D�u�r��on�	P�7�����<�,�����hؘ��w��7g��?�p������4N���������~����W�
[bOe���c���;}�������1�"�1IM��w!�����o�D^�j�{��V��Y�2�cl`�t��x����4��������L�j���n�&��>�_-]Ms0ϗ���'��t�Fpt^CHO����P0�'?	�>+{77b{�p�_{�ɖK.���7b;��R���Kft.K�&����χ��6�9��V���ϟB�3���t��Έ�E�N�����Q�{�n���Ҵ��A��S/���m������<�����&v�W��1T;�o�a(j������)��b�Q-P�&q?�w���łI�������3��jH�������y�����'ޖ�%|Cell-����l%����qԆ��o��-����BF�Mu���Im��
������ʄ����o:z�n�������Z/U�:9��c��Ag؈l9]���D�~(Ԫ����Q[�r�vs�Q�0%O��ȼR��z��M�'މ��(�:37��qM�i	�o{	^)�	�X�-
�^XU�u����#�y%��*̵3�� H��%��(�|�K9h�_�lr�	Y���橮�� �Ƅ��hQ1��g�{.�}����䢂�7��uM÷�m�=�7q����*�� iȸ3M�	>��TR����Y��
sp �w?���\�R>����3E�$�K�
k�W�^�E^SXN�|�џ(��Ts���iQݹE�i�nP���m`�RXֹ��:FW�攝s��,��X�g��v��x�<t�*z	�-��UJA,�����.��1�H,&a@������,I=������Ҹ.�ۻ���������p��w����[�6dBۯ���w}�B�?س%I�b�~k���h��<���M�FC+�8ro��8#�a��&
�E�">��7�b�[&N�Z.���s���X��<�QӜ�r����'�	�w���W���rf�F~��0��F��Fmw7!RBa���tN���VVV#�1�A�]""BB�z�֗��!i����8�d(�鿣]���X�x�<<n3;��)��{��c�q��aI���]�W������C�Ғ�Sp�&�k�l��r�Sy�oR����Es/D�Fk����kt�!)Q��zab��ކ�'q���ib��W�EQv�!|�ה2�0{zGL�?�Շ'���;Dso�/4���Q��Y�z��z*��̏�QXLX�]�tim��$�k�q��'��nO���<Uh���7�55�5xB�ݶ!(+++z4jt��$����y�q���+)���������f�~�|P��۽N���1l��[��y;�@��y۟Hg>VO��d���q9��xUQ���}p�@�_>cu�p �׷"���,�h��-�n I��9�j�FӷՂ���V�)���S2aߋ�%7���^C6<��v�y]{`	�3�I �]��?<�A'��oW�0�0b��Y�n�k+ⷛ��O7�z4L1�
���6�7��{-Byt�]�t�kk_@@��+k�.�#��(�O����+�L18������P���Zq=���^O�s{��~7�s���5���b��ЇbLXRl�D��u�N�Ţ�{t�V�1���Fc�9l�=t���9on眤�1C:I�ҙ���`�q�O��n�"�-��P��6��
��Lott����+7�X�����B�\.�(���*�>�^�K��N�v�Wo^~Uܪk�Y`��p[�V[��\>����4���@S�k#S�4@�PU��E�%�����C�'��"��y�� ��3Zhի��$C�X�n�oG@X8���g�E��v:�c��~7�;b�G����Q��A�
���T�^墡ޑ�g�*��pc"[���B5MJ̏�R�Y�i�c���=��[�?��of	��m��7Fr1 ���F1�C����B:ч0��$��h8	�����ʋ�~�?�߸q͇"�rum���}JҴ�jWS)Dt�����߇�j��;�w.)���}$�5FP8�1�ȋ�p��t�{��?��^~�eCTz�ԩcǎ5���>�����{�w�Á�G4*^H1���;>��C��33O��i��������?�������h��I�p`"@CU# R/גAUSPB�")dUS����8�U�x��54�J#��taQl)WE���jy�T�������~zueuc{�,�n�˥O�ė~{{T�
���cm�\�(k�رc'N�(��%I�e�/��_i�ڧO��֮�<p�6Y���h4�;V��;���O\�zevv�ĉ"������;t�P��\[[KӴ�����#?4�|�b�6��'< �ij�)��X ��D>�,�������k���b�<������M�
�H�8�ncp��C��
�bzd�p��I�@,�d>5"Zk�}xM��Ç�>r4/�{w�1���"��9Mӭ���y ���|�z$ �~8�*@�2F�>l����*����9W���7�,�N9�Z$��O�j6�O���ݸ~���p�$Ƙ�9�"�\v����ڇ����Ky��J��i�W�2�^ �Z� u�*;e�''�T,[zH�i:z�
��s�޽S�Μ9{���w��_��W.]>��ѓ�:����pmm�9�viz��G�N���?t��G��|�~����� @�G��$��J�%���G��O.  �03��� @���������?Z��+*�b�� ��3�!�I���S'S�IjG����_�����[o�a���*�̍����^�ci5<��^gsc�w�q�[YY���F�<	h�M��c7���&T	L"
>hs�����������7����� Q_�ƍ����W<�X���X��ؐab���F�Y��Q��
L��&X!j,,�#KN�ڝx�VŃP���d[տ""��e�����+D����B���uV���{��D��'wU]��R���D�tVA�(�FU�T�H *���XrSu� c�'@b��b8�8r�@���J_�[
Z�#�C� �̂*ƣ.� �x��:ucӚȇ�ʩ�m=���Ľ��9��٠�'�@l�jqBUG�13:�@k]�E�\��Y�֝:p!ij��SR�TZ�O �l}_��FU��|�� ��u�ACI]-��(r��7�E��{����v����}��V�V�ݝ�|V�?�2����f�� ��e�f�����ٲ(�9K��L�D�,�~@�κÇ=zt~n>p Ѧ����ѣG�?���������^�hE�����(D@ư�s?��r�X�����������뿼v�V���i��a L>g��"��}c+���]Mk��cj7Ql	��1A��΃T_�jY
��9� �Jޗ��`���3�1:�.��%iBD֒>W��<������H�l4}�]�Z�V{����c����?�j�7��O�<����u_�����vvv��\�r��ݻ�N��'�f�F��v΅�/^�t��G׮}0��[R⒇����/�sDBY�����GJ���j+\�
Hݶ}z�
J����J/x�'�jk��Nk�*�4Mz�*舱dR���U,-�eƘIA<���%�#7��hx���|�ٳg�5�͍͍͍�x��ia�ˢ�j��J�����R}�(��R���������ij��Tϝ;��)�G���5�}�����~�w_����������㽽���%qI>/r4hD�
y�&BQZ�8}M�\�q4M��x*����?��V�'e10<�/`T�,�<�^���_��_x�K_����er�h00�䩫O�<q�e���n�ann���Υ���7����ֶ�6._�|��ECH!����E!�`�D�_ݖ��A�ٙEP���9�����l2ˢD��166��,�	�4&��n��' ���k/����wޮxju��ò�EQEnCKˋ,a<�G�bPc[�f{���˞���Aw8A�������}�zP2%��������!&D8v~!���?Xy��ZKJ
H#&��Lr(��nݡVkU;l�W9YW:���G�[�&��|���g�r��J S��7�3^}��7S�j�!�s�$YꯓI���ݫ}M����Dt|���
�6B������L�H+�r��bQiPǎp� (�i�y>�8�u���<�za�Q @T�U-Ӑ�V���(z+ �^�G�7�����BDu����A����=)k�Q�_S3H���ǽ�s�X4LO�T�^�i��M�R��FE���n<f�> ��@�XD��Q>���}(���h}m}��!@���I������sDH�h4��"��!$i2��8M����,k4�,;y�����C������9�B��sι4��and0&�)�c���"��5I�%�v�����G?�˿�εk��4k4*άC��#�����:h������\�2�_P`}"�A�L�����̜$�h0��Wɤ4u�F&"E�J�1D֘4˚�0kAYc�2���/mmo�����޽�7>�����f���O�v.���I�̴�Y��y1�~��\]]]����ҠQ97�8����,%��>�#!�)K�ȹ�q�8�������U�?��ǔ+�z��8 ̕ "�����v�qĊ�n�)��b������Ӑ�Yˇ�ݔڋ|�OKu����$�10�y~�֝/�K���g766�ܹ���V�X_Y}����yb 2Tx�X�if��ťPz��&�^@���,K4�!��dQI��,D!�3�O����/�����v�%n~~��������}�������8�qD���K�l����������V�I�|��q@�zXֿ�Z�W��C����3S˛5�\̒$B��믿���K�N;&����}9����p��̡7�>0�f:��mt:� l�9~�(�ؒĘv���Gݾu۹�� ־B���"��%���$.�	��`�eJI�  .q��%P��V۵�.���W_����w�y;/
�,βl0i�#�P��e�5����Ç������`4R�j8	X��ƍk���`80�2(�"�Z�!��5�f"ň}(�1���x\���ʰ�]��e�Dh�/��e���PD�2��{Q�E"�Re��9�?qs�_�hW��s��,��PT����FL=���Za%��1Gs"�1�%K�W9U��7*�GH!F6�*~�ʟ ��a0�`�k�,�R������P� V", `��؇ ֑0z�u+̌�ٲ���d�=�5�PH�qA4� P����"i`2�FeK���Uj�|T�#5�X��N��"��b��#�(`)U\�طJtcDPw!:�~Y�MC����%��ܜ��E����p  ��N������@Dpα�h<Td�Y�5>�r+1x�d��R��;�4G��,Km%�.C�,��n�Ν;�~nn���/MӅ����<`�y6͊�DC��h
� 0�	��{F�V�����/�������ׯ�s.��Z���S%4 &Ld�<v�~�����]j/��Q�FDH �UaB�!x�͂h�4U�j$2��x�ד�(��pX���/�s�����[�/\8z��o�������HD<8|�ГO<y�رW^y�ƍǎK]r����p�!���w�t:�V�5�FFDeY�!�,�.�yd���h�0�P��QS���m�e Bc��0��D�[���KOs"���M��Ĺ���Z�8�LT��}O��&"�U�	8�ZoB�T���d��?C����>�[��TYp�4��������|���?�����8p�^�����˗��[�n[����ѿ����lo?��gN�~��7������_z���K���ڭ۷g�m"� �������g>���?����vQ�׮��Ϳj5����w777/]��ˉ������W����{����/~�</�%x�=Bz≫�~���C�V��Z@  S#y��&ʊV�0��&�t�"������Ǐ'"����e�������k�f#�$q�d���՗^�>>r8M�|���uEĹd49k�5�%��h4��a�{ﬅ��E�}��^�$�H�e 0��$���
K�ʫ/��?�oo��:&�iO��`B��Ԥ	���(}933CDڇ=��$M�1 k��e�E��������5�:&�t����u�Z�P��E���f3���\zE����h �x4΋��\l��US��/��y�ND�M~�8��G\���V/EP�q�z)
ܠ�YÓ�g����Z3�X�qB�5 ���m����()UtX��"Dk��2���BDS��Cd,�%:b�����X"��X2#f_��+�@���Ĺ$qU�3��p5�>U�MD�j��+�NLje4!D�"f���Hz��|�v��A��  2�b������H��
u|,���f}�.���z#J��)�kh��U�V=�������7��}��cl��F�����3g�|�O5[-M$7o�|睷ww;I�5H�d�~��ֳ�cDj��1h�*71��A��h�Z����8眵Z���,�BY�y8nomYkggg�F#mk �䉓.^p.��9v��l�󑖓���s���"��ڇyQ>������$I�u�L/A��p����0V��;'G��w���]�i����6��o���ҫ�!#T���K�#U�{���ADc,x/Ux  �ZM�������n�S��߻�_��쳟���>��3B������Yfy��Ͽ�ʫ�N���[jb]��<�<�A`{{���5�X!c$p�Hxh��CDI�ި���M���DL���"��&�>���>з�"�,���?���5�f�u:Y,<!UiJ��3#y�U5�e��0!m�#�'iB���:J�=s�B,B�f�'��$�?s ����p�`e��}i<mmm�iF�ׯ_����/�����Gd��>�ٳgμ������?������������ֳg���Wgk{���u��z�ݽ{��_��������?�EY�fsaq��7x��A^333�FS٧���������3�~�V�Qy��H�l6���������������{�a쿂��D��BD�9���y_�"��&�Q4�b=�0x˳UPڭF��x4��(5VD�(�,��sg���oc�_���/��O�>��/\������2/(B��y�����,��'���5��:�����E����aDh�1dv�����������޻h���)C0�~�K_�_X,��gBW�\!g���㵵�ݝ��8����e��h8�޽3�Pe4B�!U/4�M'$"c�����x����b$�L�Aga_�Dh�c֑��@Ĩ8A�K�C�GP�����&�+��$ާT���c*oߨ�s8I��3g�[�+?��(�����j�����T���J֌���RD�y�f0"hY��
��MQH��8�1����xNXu��J�K5��">Ei�!c-�53�����is��2H��	q*�5��OW�uS�m�;�����S�f�ADPD�!,=���	FĘSVj�H�������փ�R���O���NDB�YzxNPL���j)GGU�����k�|�Q ,bR ��vvvv;���m�e�Յ7��M$1n�ZgΞ�Ҵ���8��#cl�ј�����@۷������ p��^7H�v��nWK9r��ե��[�n}t�#�W�3.M�V�9;�xءc,�䆣��~��^x���;g�Ě�����*���.��=<1ә�h��,��?�E�ՠ%M�{�^j��΄D��!���3[ksQ�e_ۋ�(;>�sI�ć��nmm9z�Y[%if�VVV���Ed��!���E��䜳�j±a��ыf���݊y8�ϖ}i���DqG:ȭ���47�p"u��/�3U6�z������Ӯ�e
@�eq�*G�ʃB�""��qH�9�0� _�^#uQ�Od��X-F�TN(\����GI��<ϓ$}�w�;v����C��,ʲ(����'�f��'�l��A��eo������������~�[������ܽ{w~~�����[��^��&C��D�W���?������+���`08{�l�f�v����Ξ9{����W.��=`����w�����yc�ȑCO\��l6����χ�x��v�������;Y�i$VQ)j%B��~�Ф��G�S<�+�, kՂ�فK��H�YD)˲��Z��KɲF�� �؀��������_}��;wo��W�������u?��~�&Κf6�u��l&B?(��tR^�����������V��U�������G�Ld���^|�W���|P���JeYyq���~�ke�?����%#"���;z���V�Vo޼��I�������
_j6�(GAŉbOTE��Q;�D,ˢ��<���T�n�X��[$���jZ� <�5�,����
���I�3K�~�~���$"D�!�L��Sl�Q�L�W�jzv @��'Nm��,��d�H`T�8�PU���������Nr�`t��"!���b�Ê>��@����%��ƣn ���È��d��b$��S�A��Ds�yw��T�1$�B麥��V���Z��m�����"�)ϲ>N%kTIk{�Lj��Z"*!T����6�P�{1 CJ�G=�t�Wyv�j��®����LWɊh�uѐD�	C0X�uuChL@o "�d��v^x�����ǏYUX(�uY�>[F@A��'N���������7�������s_�◾�_x��?�î���v���,��{8PI�s.q.�2km��k�Z�/_~�g���/
K����ٹ}�v�Ֆ�|$i*"�о�F  ����{_����(O���j�4._��[�KKO�V���|��q�ى�Y��c?Eb�>�J1��� ����������"0��q�_ʘDc�E����/˲,�3����:�B�����++��d\x�� >D�26d�s1�E $�	�K_b��E,�09�f�d4�~�r�N��}�Ak����T�.��<V
s��Iն X���멸N-�>�b�UB$�+M�8�Y!�<E:Gk��������DQT�,p���^b�q��#��-�!�������sEQ�{w��ş��x�g�e��a�����������B�k�w���Lѯ�������"/n޼�������`����!FV��Ͽ�����G�K�����������]������ׯ_���WWW|���������sd���^��t�9b����������!"k�B�z�L�H�CL6n�<�ۣ�qܞ��x�?標�2���v �j	�K�9��|4�www���N�:}��-"�ƶZ͢($DR���hh�����X�r|����q��C��< U�q�L!m�oc}"��!f~�ͷ�����q/�R@�$�~��/�K I�ԗ�x4ZXX8�����#"�._>�|����;|x���۷:�N�4uI��Ď�1�OJf怂��ц�!�L���>�ē��3�n�Z[[!Ăw�,�Ν8[2߽{7��ھ�>��B$B��mWT����/�
�`ʂ�5�LC"UrWߨ~�'o�dߪ8]�0x����G�Q�N @�jG[�����k��~ʲ�Z����^@@j;�@�$V�Kj��F����?S49��HD�@��������caCbX�V-�!c&�GWW-Y��JiHAKO�1 Z��Zy ,�[_8A�b�x�8 1V ��
ԛ���f�	�1�⃇��T%���R9_AHU6u߰ �!���'V�Tb��Ӏ��w~4S�3�D�d�780;紗q<������^��N�	bk�N �2*�HH.�Y#C�T-�Xg�F���x���7nxDF$�#f^e�����U�̇�!6��N������l�"����n߾[e��s�sssYc˒��d�����u��E	E@�D!
U�ǭU[��)��uS��V�3&�O��� ���+㹥��["cL��+u�M�$I��,��Q	4x N�����9r�y�e���*$>�e�ACD�4l��)zϪ��!h�[c��H����D@]����"��ք�����V�#0DG�r�4M�VLy��"���8� !�Xm� H�&�tܯ�PÏ���O���f�H��j�^,N��1�,!"�l��P�c��p\�+���\��=�*-<ST�C�A����5.q�@��A#���;������^��\�a����:�VK�:��[o����C��$Yj������4IѠ/K���1D�f�D�N����h�>��(�"��G�_���I�h8"�����;�+�eQ�i��˯���[,������^OX���"��ʢL�.D�JU5�b��.'L�	�F0�CN�
JN�깩��=����u�ཱི�� �d�4��[��O^���������X��W�2�c?�2O�TϾ4MCB���/�_�L���z�DY��l"��%>ȁ�0"L3��An���S��Ngw}} �4�F���e9���޷��gN���*�d�M��c-�żj�
p]�
X�eQ�f�[����>�'��O���J_*-�,˹���o���������&�"%@���HF-����1~FU��l�Dhau����Ӏ`$-�(f��z&^]5���w���o�a�s��T�G���IE������:Ҥ=L�g՟ ���(�'6h2TƂ6����1*�U��h��K����0T� ���`��b��bFf�+��v�	�y�����
�V�B̪��B&�d}A�&���U�	�]E��!V�' p%]�G�r��-
gL�R�C�5D���S�'Q�"�H]9�~�D�QD�����x�Ax(������`TV�~c�� �,KT�"���r�����_�k��Z__#kt�]��W__������L[��s�,< �1%C�TDd����C�'������Ng�����������-//�+_^XX�{���ܜ����e	�z�"P���[g�1I�m4W��pј�k���'q��G�U�j\�j3�D{�H�S5���O�B4R$LIN/b`a����:c��5�V+�	�Z�km��yQ�Ɣ�5�D���j��[e�*lDDCG�����(��YQ`@���32�h
^뜣}����X�BmH'��~�R���!xo����F�~e�#�E�F�4Tݷ��y�s6=��F�" �S���zW�{�&��S�7C�:bP
��r��E��
R��c}Będ�+d��G	q����W���Y�i�5TӉ��V��Ȅ���?��"Xk���L����"��6;�,�J�x�±��ĕ�$g�!Z�[�[@"0Ʃ8F�/K 0�q2(�~/�l�t�*�7��(���hTy<R�6ʫ! ���C$i�`�4H��	}Txb=q��d-�J�R}�V�y�y��3�Y�3SSå� ���!s�������ǎ�cD�s��`0�9B 6D�}��g̸(�٧_-"�9f�tF�@���@�^�dC��/�R����X��]���%�EY����9"V��("���/�<����������Zm�|�&���4�Ԓf0F�5���.�V�bͶ�җ�"��jM$��}�| �r}S���Yb<���[t��3�:*�����O/-�S'�,OǇyw��S>4���ea��:[!�2���/\����C( �5:� -"��ۀ���>m`=����l�E�Xc�T@+H"
�uuq��ѳ$"A�iz�z�A&5�qd��G�ƾ���^*��T��5��|�kNA�>��#�6�>�	� �hC�����#_���(D�D7E���V�Ru�����RG�j��O��
kE�+M��x́I�� R�'�"�����z�7��n��,F1�eQ޹}�޽��fsvvV ���rQ�Q�ܐz�j���`0Ȳ��������� =v�3��̓O>����������$��p`�p�*N�#�&I�h�mBt�jJ�z�5=Ac庑��ձ*���*)�'#2FS���ڽ���i�̾��"��j\��K_r��rEw0�� V����!����4M�/}��d�YD�o��`��0 �c�>��S�|leF�8���H�pE�֣�/S�U`���ODHDB�߶�qjT�b�֞"� K�z�$�X������8`FD@��(N}�7�c�k0��Q�Xk�3Ab�w�j17��+��נ�=E���kL�U��\�$�!����Oof�\}��KW��8�T*cd�0��}9���>q�K�x4� ��s�f�,|Q$\1	��l&�d	�.��` �"�=�U�j���%�EQk�ebj����N}m�U�Pd_r������'L�]���e�P���Q~A 0���6�4��^+� B�����*��%�6�cM4��"J�D�LG�*�x�X�ȕ�ƧR���&:��*� h42RWK�i���ݓ3E�B������PQ<#1�P���s�F�����~��w�����p��o��Xc�2GB_�EQ B���D��bY$��ie�5�
�~�÷�~geeE-��cM����?�2fmmMװ��XtnX��>��Q����cG������5l,�N?���:���U�Ժ�$�l���7�K�=Gi��^��Z@�3UF*:�?� S�\�Wr����á��Ȳ��d2�̂,���g"R�z.WLD�*�bTi�3��$�d�9��[�$@Ԍ��NfV�&T�r#`��Y�G��o��׶ TmJV�>��cNa�\�s��S���P! z��vQ%��q�p ��,4u
֖�Bε�De8�lBփ��,P�rtA��Tx80{_Dͼz���ԥ��"�C��s�J�X���� c@���<k ����'��r����P�šC��4m6������������h4�4��&4S���NCH*=V!D���U!JT��xN�ǭ��ZKW� ��c.E�=|�#uj��nǼ(F��x<�����!4�=���k_��y1������`�~�ȺT�
����D�-�
P$2�F �xq�hRR�<R01�ڪ��T�~����'�>DD�s �d���o��M���h�u����Èm��R�n��y�#]*P�1n��WE�KC\�:���
 ���ܟ>ّ�������
$�Hl���*�H���ͦHj�n=���4�����|Ҙ�왍�~=3Rol�M��\�X�ZQ�L ��-"���?�D�\P [z6�lT"qoĉ���s������(:%N閷ЛN��h��
Я�4
�OZVec�0�����HV��ǢiD	l>�w�� s �ʪb�5�D����!�s�AӫE����o|�P>�|��.v�	�<Y�\��[��tfDG�������($d����R�6�A��MU��ƥ����Ĥ�4F�Jv b�B�P�X�k3a]2�S����b6��O�t��#+�������e,��C�C,.^z㫼�y<����dچֲ릳�����[7��"Y��� �y#�qVf�1���փ�ؤT���ܶ�G�rX�N��J�[��1�N��@Dŏ�
 �Y)��w�3[U�IjO�4G����6H[M�o�n�6�ќL%�t��5�J�;�H�L�A�h��I��Dm5b��+
� i�dS
XD�����̒��
�UA�,
#���OoX�)�n	��vc��M8B��b&��cm!:�Q[���ҧ�"r��|Z��
`Dꐈ~��2`+�jY�i~%j��<����K��m�\��� ����O�*�e�>�HA��q��Nʎ/s���<��k�sD*8�F�H�n� "mB��l��ɨ,K;��)7�V��(KD�ED`ns��Ԋ�E�Ҝݪ�D�;wvm���*1����L��m9�� �Uo�!otk��{`�zΙDR��x��Wq�8)�
�43�h��7��?w�'"R�>`'����9�=�Ʃl�����
�������sq�s�.��R��A���,˲�ȁ����(��m�
�:���#vy_��*F�"ڝ�Q��[2� ���%� ����e�����9g����
.	���2�i�pD�����C��bm&Ċ�6${��2:�8��y�NgTH��*�Ћ�D=�t2��!bዦ�Y�棙G�J ��HC�q��ãnU��HE9��d�>�����.�C�G-
P�J�f8wr#c�N��an�	��#�Γ�4� �#�Y�	�A$���.���NLª3���ɵ\��p;���W�!����0��1o�д�b�!"�rP�#��&��Z=�@�9(��i~V^F�  %�I@�Q�#/�Й��n��\
�(�3&;!�����yd0j�l_t3���n�Ⱥ#�0	\���8����u@T��s�����ht("�n�@k#����
��<8�
H��l6�$���e����LQAQa�җ���J�T�Y��4��cc�v�����c�c�x�{�Ǜ�ߕ���r�R�a�IU����Xn���ǭ�h���Hnf���qez�ƀ�t]�;���㔃�$�C�R@�3�تљU�+B��0樠!i��9h�(�<��ԥ3'�t&"Br�{_:#�4�Lbw�>�2X�C�RR���Q���7EV2&�L*�(*
��1 ��3|+�i�@����D�%u�� @�h�cV4C@h�\"L$���ZUEQ���MӈHUV�(Ǚ��IQ�`�L��_�/mO�H��u�oi(Gg�%F�WX�&h���i˲������ ���EY��۳��U�\S�ׯ_o��ҥK�*����;���p����V��kg�:�u=!Te����9�����Vn�i�
m0�!a[�
����4�j;ٷ�m� ����!��E*ꈻmο4�*���>��
��qcD���D�|����`�$�	U�p���la0#��Z�໥��P�=�K�K�t 
�Ô�,��h�2�)BRRIPR�����C<� ��&_2&{�x�7�e^�H6a#��R�������"�eL�����L��E� $q���A5���  ��Ų�#�|t$��g�U�-���vm��1��ouE�JTɋZ&��!�<�#"1�� ��0ř�7�G+�Q'W1G��(s;�>? �>�����UP�!;�X�q�H�z w�e��U1$�%�0�Y�)�/�9۔G�`@Be�#�j @<))�*�pc޲U����"l��HxD���Fo  ,x
B�X��[d��}�s
Z(�M3O`kk����d�"��hooggg�n�$�����y�@K5@,�@�����4*��"�yڮ�?#:UTVn�PQYP�!�US�����M�u�F"!�,"��Y2�R��gʋ��y��e�r�f�Jq��!����2crq�s���|`Ml�6������	��ԇ��$���#\1O=����Z�{_�%�6��%��n>����5(��>��AcK��$�fe$<��f tΓs򕔖���;v��ָ��7�`������'�,B���@C�0i�tY'rP;k�18* ��4{�Å�`�����kkk����萜+ʲ	����p0��W�r��Ŷm�~������������jP�o�����4M���aV="� 1�z�����H"
��Wʲ\XX�(��Tő3-yTC&X��UQ��y��cmۮ^A#૪j~�Ŭwvv������ʲZ[;��3�,..=|����{���ZQ+++�Ѵ(�d2����?��M��F��
MK.��P�s�,u "u�}�YQ�v)�s{/�-�c;0*����ǦXc�3���R��HQE��3�ȍ�8%@L��"X�Y�bMM�!@��^AL����yiDK���Y���?���s�y#9���e ����X���{'��%YՏMEx܅}���H���Q1�c_v�N&�m"C�t&b��Y���������LE�O!���Q�d>�,X̦Yo�a�˲��\��5��#�%OVځ=+$j��=���vp94&��˲,��m۶m˲<u�oh4}�[���Q��,9�2:y�G~�I��Z�hY ���w��Z�|������P�ɣ΢� ��La�k��)劥-z\e����["[\,_Mo�9���;R���<=�ͷ���y Z!N�H���[C��π�+E+^H���z�Y�sh���?��Ӄ�������������ht8����ղ*'��	K���0K��4�
І�4MUUf˚�.,�y�ش��T!q�XD8���^�T5W�j�Xu�����ie#��8� �jf��*�eҞ<��tz�r1)�\�O,�9s����8�	��-�B
�������6�,��ꛩ�cxЇTT���xO�<��5��?�a��{I�"D���K,��%B����# 𖠨?�|P�� �(K�@I�16E!-�&@�ؖ�r=\tQ���WR�� D�-}U�E�|@$T6���	�D~�8�s��Å��_~ّ�w���O=���O7MsxxX7�(ܹw��ࠪ�g�}��g������x����v����?_�f��˃����O�S�-Ȓ��=�t���T$������,���U �N�Ӻ&PBK�υ���m\�x���E��>��۵}\7MY��<�����v��a�@F�8�&�&�i�4���8�L��ॗ�����_}�M�կ~y������p8$��a�Z�N����˚^Y^y�ʕ˗/eyx0��|0�ή�={����PD�_�~��=dֲ(���n��n��9V��6�T0�.�'�5�tD�)*�2."8��5�B���" �QE�lIm��~6��}Y�E�mD�jH]b PAz�D`��Q���W �X-�Jh69AlyI:G���|:�8�s(U��w3D0O]����q��~*L�[\I?���/'�����Ν[�YY���Zg�����Ʉ�,;��p8�t:m��(|̑&.�"Z�:�S.��)�)��d�4�0'��s4;��l9�M�Z�dZ/-.�e5�LV-�Eh	m�9dVh���;��<r�d"rVř o��H2b�cc��ɳ�����xzK��Ʊvޠ�'f����`��c�!�|��:/}��D����2��PA���uor�P��fsJg�w	A"Ɏ#��,�,';�V�%V�B���*C-�2�
,eY��i]Of�7o~��������+������{���?|������mYzp��Մ`�-h�Z31!��@�T����f���bAEQ�o�v<�e�R2��ґ����\�"S]����Vkj�Շ�N��;�6��U�
zZ6fOG(Ԋ���[�LU� ����� Pc�� ��Op1('���)��� ň�a"H�O���݆ 䏬��Hfv����?Fj�$�ⷀ`_7�HX#�s�����0R�H�7�	C� �^i.�'��\Ӛ�'ْ�Ǡ������6p�]��9fn���0�V��a���d�+�
u�x_�={VUWVW��7.^|뭷Ǉ���7{{{"�Cĵ�����[�n�����x<��q��7���ڵ����hd��e��	�'���֟@�c����	ATb�iG��C[܋/�����_&��Ç<�*��Jή��������/���g7o~B r���*�o#��D迼��06M3�N�����ξ���_}��w�y'��p8��ݝ�fK�K���Γ��Oq
�ʨNɄ���ٯ}��ϝ���]Y]������ʙ3o~�����u��z�������i.]�|��������-����{<�յwE�ۀ9��t򅱗�a����ُY��驮ts1��y�'�9�l�4��RB��m��/ʒ�ˢ,K�"���ղ�	�9p"�C�����,�(��B�Z:�<�q�
2Y-��bNΗ��3,a,���!���6P���@���:�t��E�e�(@�Z��x<Z]]��`�43��ϙ����S"bDX�EY�u]f��b"m��D�aP��UT[@�5��hq�8ť�%@p�;
��P��[pw(P��C�P�h�C��w�1���̽����$sb�>��g��c���c1��_�n}@�u�/��X���Ѩ �+>�Ov�ţ���������62�(��X�����cn�Y"n���or�HiyH�t��q<��T�Ξ���-+V�T�������I���nM.J��崜1��kכ\��=s���I�oK b=�MqE��C|y;�t6�J�k�k�r�I���������,��"���}���BB�,���]8�	��Lㇶϼc�t'��N��"^�õG�PY[��@{DL���K��\��q�[�:�׹���^=���c�����a;Ɖ�� ͂6����?Lt+!e+��aLLbQ�0&�f�y�/o'�C�/�O��ks�N�1����S��(���*��`?39un�@��4���; )��=P��<���h䩎���o~���ͻ9�'{��C��9����W��_������z��V� ��[�3� �w}]<ƴ,�.V�+&O7A�:����+�+Z��z��$���U���y�m�}9 ���R��Xҙ�05P�577�9����K��������n�}#H*Y��l��"�G�
nnl��0��M��9St��!7�E!G�	�����y���(&&�Ԁ(+�D�����u��}�@�|�P&<�HW(�Ϛ�.dA���{p���w9����q7�*ssxT��ɝiok��ME�Ǽtbp��43���J^z�I�^k��oK������қʮ�=��P�2js=][������>kvX��m��a)G���NS�Vz��ڜ��D�g_V ���"�`�y@!1�������ȝ?K��*$6ʡ �0[`ЬQZmi<P��Ym)�Q������5{��nu5p���\��d��'uH�X+nw��#�>ҝPH�2��>&g�oGH��ɴ�b��Q��͋�Q�ˎ�Y�������e��(h|����KCiU��#�Fb�'��*�[��9'FZ�w�+�[���^3c�L�e*@�7iD 8N�ዑ��7N�9��$�{l��o_��$�ۭ���4;� ?C��)�!�>�JYV��2�:| �XO	Σ3��@i>�E6J��� ���Z �w]c
����X	�z�E.?N��e��ݽ�2S��H������ݕ&b؟�`U�O�,��)�>(h�ѡ���J�Z&�g�[�y'V�W�MS,d�8�>Zy�栫|�	���Ѓ	�����x��i��~1@(����57wv�媬�|:G�JH�,���9!�j���w3��i��N3"�uA���)g�kk��i�����d���K��O�:�&;��0��ॎ�zw�����s�ؔt�<6S�M8��Q˸��/�~�c�/���+�t���KҪ�z�>����9ԃ'ݠ�W��{@�샟U�nstg�0|H���2xd��X�+���x�1O�T��rU��k�[
�!^�Q�om|hL�L���&c�U�ҿi��8��ӑ��P�,��RU5�<	I/:i1�{8�D�����y��G��E�E>/�:��)��O���'�n�655�"��Ч�J�ajգ����c����˄�V��n�}�kO�B��W�Ѭ�FϦ_��ݺp��{�{4�&F���)Y�*�S5�f[�.���P��$uɻ�kUsgk�ea4���S�|�������c x�Ǎ���!+���&C�zN���1�W0��������(#Ul���t7�T!h``�Dqu!�2a�qy|�f��W�Iu5v�(.���h��� �
9�Hia�<�>Y]]M��d~����`]7��{]�\�ll���/!���Ʈ��Khqc#�=�-�r ����9B�IQ��2�1���鈠�ӈ��?�)|��mNWX�äXzi�G�ȡ�ZPb_6�z<N�q4u`�i��_C�7��Bs!�;�w��>��&�p���b�un@!٬��0�R[��=ؐ�4c�zr���ߌ�6KpJ��zN''IE辒�/g������ Uy\�-�t�V�	|A]4>i�K��Z��̏�ݔ�ǭ�|:�?��aɤ@T=�՗�pXfj�;%;W6�P��ZJ',U�P��O�V����+R9ý�Iv��=.��gg������<C�3T�٪`����s�㧎�*�,2��Lu��V���N�qi��~tk��Z"s�W'V� z$���w�LZ>�e���.��ۛ���b����!��Ss���M�}S*Ԓ��s$O�!%���]~`��a�K�5�zUPn��NE�8��i/"�ũ��\����d�������Q���TA�:�0H-��Z�*E[��<�`d)4�)�R�$�9��{�,3]k��96Ĕ�K����v�MiR�ʞF�<���OP�����7�5uo~^"B��f?(J����	��Ǳ�c�"��j���v����;�j���1�/I����a;Y���*@
��7�#7�n�YD��ZA�ݓ6P�h��8|5Э5�����:�`���¢-'p'l��>w+��i	X[�q%`���g�;��� �z�Q��t�F���O�+ɳbJc����z��[Դ�#�N�Ep���>_-�=��+��:d�wqvvrr~�s���_W__C@΅�*Y������܁� �Di�f���K����J�Cݿ�yf�L���Z�k��M�.�l�R��q��ZWÔ̶]u�t�?��>�0
�c�t8
v��g�T���X�g���B����4I ���4Qr��s�y�����ߍ�:��Kا�/��/K��u�ߤ�����0�{�򩬃%����t����L�Ɉ�aN�Q�����Mta�3r/୴�S�����D;,��)5pp��dM�L����$Ai��Vϥɚ�q��x¤��E�4 v�� �JR�Dl'~�u�d�p=�^%���,�[Y��q�^»�
�����V��U�5=<G5��M܁(�u�ۊ![!Z�H�_jU�Rx��"�5o�~E��H&}x*HA�c>#<�*k��.�_'�x���a���f ɽ _�k���4a�i����JN+-�AʹK����9i�k��Y/�_�7��ǜ��@^�ٷ���[0��>����PQ�"��Z�j��q`"����C��9��d+-5G���"x����UdxXˀ�R�D���lS��C��� ��L�Pk�J����P�`��I_��4Y�V~�N7�<V���Ң��X�V%�� Z-�p�{CE�Z�}RD�iu�]���o��j�-4��V�.���M��c��^U	�_)
d�#�'O����y�f�_  ���O
D�b��4p�t[��m٩�W[h�"z8;jV[�����`l���S�t�.��g���4�J����<>=_	���؄�}�Q�����5%U�*'O��x�����,gs�oS_��z#����u.�6]��O��
���.��mꂗA�{î�ʽ���qp����Zxw\�����a��&=ᔷ���LַV;o;d��'R5]����X\s|�J���o�n(���3�y��B$��e��� AQ$��54sYUn'�������Q!�>�]
�Z� Iq��7������S�EG��Ôg���_����� %�%i�{�Ͽ�Y���J��/d4��b��o=�����^ ��MhwU-�q�V��	�>��"dAwCW�M�x��]3
�������R�)ԸF���=�!�EȼBmq�l��PAŌ��e��yPɘ����sx�GNZ��֥bG��QW���`>�A&�6`o;�n/�sMpi��'9�oIp�V��˻]d�La��2��!�K#'#{����u�����abb~2���jq:�)׸?Ԗ�Z���}`����-�r���y�0cp0�����z!��bDn�@u�ęwWc�ܗEg��ݪ\��f��Q�XbWч=�äi>�+]:�D9
<�+�_��YH�TS�ͽ�M52����@칃6��5]�Bm�n�tmuĢ�-�b�-��/���[M,lj��cӐ��Ƹ�ّ+����d��"W�â���r�t���}?���wū[r���o�;�=7�����VV��{Wz9$�����,�nm<�*M�Xlw�_յ�x��Ӻ�!PDF��Ѣϖ&��(��o�2��]:.�C��9��ɏ���)L�����la����Ǐ�`��3ܷ����ܜ�:(���>a�TW���h1 ���9�0Ɣ����Mh8:�*����z�ߚ����^�M�v�4Gd_K Kv����4ɑj�,(�Sh�:⡕j���Z�����i���A�\P�e��д��F��Z`uV�\v��������ah*D]��8v���EH�wr�Z��<{���')��q��ъ�dZ����9�K��[�kXr�]/<��C���4|I='�� ���"�Xd?���Ol?#8�$�ai&~g˕����r�x��<D'��/H�9���L*�9��q=꺁k�~q�*C���Ka�
����2��ȟ���T���[��s��=��;>d�&3�|4	umQ��+2&!��F�	y#����Hm�	��շ�R7�ϵE�m�^eM�o k�F���n<��l��z�E����h����ԏlc�~Α\����6x�d�-)����)��|A.��$]=�%���G���ql5T_ږi������M��C^��π^�c������ʖ����o�1a���ԡ���S;�Y�݋��=����ߜ�ߠA�e\�O�w�;ͩ����ΦT�q�vp�?^cҽ�����A�Ux��~�m�i�;�:�BY&�g��[��%gn:��*�_�C��j[��??��D�y=
�
�Q�KB,����8�;9AUNI�Y��4"��C�9��?��j���$�������p�5��/7;,��sbm�.྽=���2Th�����F�Q�W�R��`���$ʁU�b�h����S2��jք�����H�]w�@DYv���&��ب�$��n_���
椨ev��Z�*y��ѐ�F�h+(l�Q7+���sU��Q�!v8)�,u?�]@�Hjq�QQ��N@��ma��Uٵ�&a�Α�� �>5�87ad�V��(S��y�qO:� E1�����D�4ߢ�PDG������j�R�-����J��&U��f�h�B���>E|1>
�cgIs�&y�*��g�Ԕ������U@�<�X�F��h@���dMm-���Rь���;mmU6k�����qF��@�CR2�v�Ϛk���2L��Kv_���\n6���[�	?�n��y_�g�^/6NI�I>lb�=X��B���m�L�J8��4�o�.�i��\��&�'�WߴKȹMM��.]����F���?B_��/a�0*�E+//;���%��맽=W���6Jϛ//��bT࢐ rd�.//7~2�BE���C�1o��{�s��x-���ꁐtl��ON�Ul�Q�"Ë\�y(¾O�!�����Z43���4��R�H�������e�h��i�A�bI�0�����,����1Gm�������f1�M�qL��gs�Uf%B�N���j �I��,p�Ղ�%�D����M�(1�^�����΂�7]l�|{�n����3��sf��!JC!6�'�4�d =G�ܿ���X�_Uh�nj/0'��U�i:k�9�^�Ii��,l��Ff"�*��i}������(EZ�A��t��y,���v]3��_Q�/��Ѷ�X��F���3�oG�q� J�[�����t4Wx���F��C��c�����$��	���wǖB���;:�q^ U��V��_�P&T&^")�4Ԁ��K��)x6ci��%a�/��Ҽݛ�,�~�d��A}��l�d5G>uuja�ݾ7֍���cܽ����H��9��300��˰�1j'
Q)������l�7�L3�L�'���!�&<���}�U2�2!�C|�Ҕ#T��)���{���\U���& ��:�������H�D��`r1������9��e�V�F(�Ҩ������R�=�.c�{x�	���NOO	"�$Ns0ޟ�פ��ݾ���b^�d`�{�_�Y��Ŭ6��:j�N���	���ss!�:��
���r�ݘk�_|��L���6����y�%���nk�)X/���Wq�ccc���iN2y�N�ײ�O�>�&9^B�����`Y�{V�
��f[=��ʸu�T�hu+�Fr��1	����t�M����vg�-�ؼ���&��A?0W)�Ф')S����d���=�͙����+?��	}1dR��C�\�:�L�*�q2�*�p�*��Ic�a+���-Kg���3SJ�sUm�{.�z[�=?}�����ρO���o�V����O1�����&FF��?KMM�st���}��.��+�� �ޮ���#$Pp�}�|��AԚ��e~��sr���S�&�5AFF�����}��DR��^ڟ�140Y���:�v��%*� F&>�WB=9�]�g[��Gx�
�7MKK{�{At��JY�<
8�7�ѯ�=�^Zu獞�Ye���1�fZ`\\�H�����|$�3������g������R�41�i�L�1��A+��s}Ќ{D���j��5�~{``����z��OY^����'������4=�ϻ�WWW�WT��.j��TK���})�i:��s���orL�8i�>���7��ɬ�X^�Ƴ�k��쿏�����m7:$H-ߢ�ov'��ڊ�r�G<z�wF���������,�O�(�-ZF']�v�j�����Ǔ�<Q��a�!;E *�D��q�DR$�_Z|m�k�K�MVO��y����5�J�X8�c�×���-���ː�i	�)t�Os^�q1��K�|Q�%P��c��:����D'N�m�_`J�b�Hb<�2���~r�c�I>6>m��	��μ:�A�-?�*(T��oI*!ٳg�4��N;��N�TpL��α���! ������̉�_��+�B���1�,�-�@>OMi-	�0VA%N���R�	ct����d�����L �
"��#�M�s�{�!���K+g�ט�����~���<g�}��|>�x윱5J��}��eW�x����˚�1���9]_v\�(QN��Et�M*�q���sXM�<�X͎g�e�W��*o�M@�^( �}q���'�M/5}���A�7��8=��b_�9�M$ɦ��|*(܊̺p�KE�� C�!��������	͔㛷����Sw1꺝C�>���������mu��}��Dɤ$� ��B�w�"�����R�Vx�XaTlT���b����I*���8?���
�;����ϟ��� ����6���3U�v2x#QJfpd"_�P'J�*�gg�[	�C��}��6��@���e�w�J>�.��B2���jy�����c�X�2�5�o����j�jU7.J܅o�����#e}�Ot�A�D�s�bb��\�i�M���Ĝ~$\�i�oE��[�d���\����N�Tc�ۏ#���ňzcհġ�_e�(���O��G��N|����c#y��J��컁هx,B�Ϛ���I�M�3�@R�oo���W#�1;گ�	[�~J~>:��G�n�o>/�x
Qs�߼��*eI�0'�������%�59�+r�#y+�F<� \�վu���������Ε<}��ZXৢ"7�;+aO��^qx>4}�4}�J�ғ�N(������^�ĸGA	��5�#\h�*��0`��^�v��SK���$~n���߭�����X�z�&6�)��^.�ҫ�j{?�/H���\�� *���_���l�]T�ZZ��m�����`≆FF�B�����j�����������$�u4}<@�Ȟ�gxI����(.R3�>YCI6�. �^-�xë����Ru9�
��WT!�P���`���,�ɗ�(�	<��g��ig,�b�@�-��{|oു�\�O��St����zv�����U��1�]'�T�H��kJNmdR��%GƂ�Rӧ�y�&h_^���,��Z͍�'�#�Ǖ��#j�ɹ �:�� �!�Xj��c�TiɚCY4��W���h|P�$��P)�-v�Oa���s�9�m"(�k����Z���&�	�l<ZD�r��⏑J�!�?N^��>h�EDb�h�A:Kp�)��}iX�:����2$���G��Y|��L�cO� gy��WA�Z�V��v`8�a��AzJ�Y�&֛b���OW�r@�-��ٕ*�z.OGI*Ek�ـ�_�����=��4����Ŕ�+�R2X®W�-��y�5X���1�@A@�:��.�v����|����76$�N���6S�v�<�q+-�FԹ��9j֓�z�[-ߛ6�e���t�κ:��c��/v�ɱ�S�`��d���=��������1��b�b�{��=k;���%C��ey�C9 ?7W��^��j��Wg?���)d!�����δ�}��N&sļ\62Ԙ[��)�0��9����E�2��;a ��m�I��82�Gkv\|�Ѱ��~�i��Rֱª��t�����91�o�#�/�8]�䪴81���d�!��c�W\n;Jr/��!Jp��� liŨP��'�@3*bM��%��N<�7���8[�֨b�~L�D%*��Shvh� ��	�#��c����<��o4��*J%�����ݱd~�\M}�GǺ���Lq޸e�%U�h�C����a�Z��U��F��W��,�D^&3��
�w��I����/�j�$��6%Q���k����K3�J���=ݪ?픤��j���!�g�Ӆi�ܗ��aV��,.<�$���&�������@��rv�$��$��Mۗ-=O�ԟ��j�Nz�$�$:���(]�3��g���&+� �^�#��y�鉵��s�CQ�]����S�hĵ�6G򡨶��yw�?>:���.%��Ј���@ u>�'�+��i+@�F�@QڄT]ݯuvGK&��kw������������J�Z��ۢ��w�I��[�T�g�v��益t-��s�5�PCCY�H��]����l�Φ�� �9�Q{���j�ͫ�<ĩ���L�����eWa#cc	�!�-`��z}[�;�F75�GOr�b͊�:Y�*s��ϼh�9�����o>i$����
g�g��R���u��7_��������.G��1		r���FG5�c
��_W�����Z���Lhi� �9K���FX�A�Q�� �����WR���TT>��
�Y\�pB$��
�r�p~U7���&'�]w�BH���z���{u��[��gĠ�������b��C�X��=� �!R�����_�n5��똰^�ݳ��#�_��zC�VY@���Z��+�D��Sb�ĳ�W�dbu�-��X���ġ�V	u��_��@lw�%y(0�:=��S�3�u"v��1u#�Vl�{y /�ȸ}}�� �|�����꽛@β��D����"ż���p¬��k[[`����"���.�{���)B�
f���e9JZ�ͩ�q�J��[�;��Y;�I�0O8Kh������9�Y�4�X�#���d��o�4c�z��T��o��t(��H�nˆ}�V6]�L�e���o��@ K�l���x^����< 恶c�	�GMty�ׯ,�`���f�[�,�ǘr�5�ru�6�J׃R��H�8����	����r��E�^�҅X�<��&��w�PAyD!��9�����dlDZ�_��T�S�e*�J�Q+�z A�p0U2���֏a/��Ayޤ1�6p�[�Ġlkh�Ax$�4��q�����kg�;�Ptu���ק�= N.1r5��!�
oEō�)"B�ڲ'�u�~���82͐�ظ!]ܥ-�u��Aj�,��� P ���y٬I��kp+��=ߺ�>�I>\�qrrJ^���q��Vs"��6�cx��\���A��%%Vr~�)z5&���7�w�y�Yk�~���$������$-;��$%R�) �o�n$o�����S	_#z��q�=�}7��\���":�z�+kՆ�ONN��깛fz^��zC����t��3��]@*b(&az�߀�v��E��q�������o��=Ӟ�@���()���0���뱹�t��YH�!�\�O�=j����������?�M��,��-�1����m�!o�܄�y�������FHH����ptԡ�G��`���$>)��mL�=t�*ݴE�Vw�j=���5GP_`���Nm����w��6u�|������>����(G�_�	�|c��ʈ����������B����T6k+b� �N���M����� �o���3L�ۗ�t�w:e�x'�򺪦*�����,�)�����g_L�fH1�(k�r�t��͊�~�k��i���3����}^g.I��\�~-����:��!S@�x1�Ą�U�jE��!�*���^s�(HQ	c�9�aV��t���Ou�Gj��y5?���VZ���� b�u��^~^�����?�d��k��7��
��D���N�Fgb�:��`��������p�MI��T��le�&^����I)�ě:�E�����nYIT(�3��w���͢�[1T�>��k�qq�����r��~���~������k����Ra����m����x�`�<�2� �� �u涉ֳؗ�/��MA�E^Mj�3��V`e}��L�*��^v��,uq�������4��岔9����!�}�'C����F�M=۝#�����#s��\�3l���躺�fx�l1��Z����`?`Ts��	�&cņ1A��CRAB���������[<XtmL�Ĭ�Č����ѩw���;--@��c�K�.����hĲo���:u�|��K���l*���z�ʲ Uh4��#�����Bw���_�A�$Xg�¡wL�|��9ةL*%�ǶK�
��<��X0U�\��m�M��`�q0;��E�������b���2������������f��﹟BE��/H��c�R�i�</5WMm-����%�_Y�3����U�itG6S�?�p��2���E�r����_�ԏ�-�x9g}�	<�4��C�r.�_�~!Y���@���Ī�D�f�/��_�󿈽�l1�SL��ፇ=�Z��=	�*G�Ӯ�SŴ#�F>��������	��̌zm�O���rT��Zk�}9ىx8��t�j�b��n��]��A�ih�	���n5N����;=E B��F��!�3�	t��(�k��:d��z�3C�/��u�R����c�9T�L��-{xy-�z<��-.�\����ln�M�wwu��g{��Ϯ�7ޜ�����J-N�k��J}��U	\����ֿ�iz�c��\d�ۯ66����0��ՠ�:�����n��>s��.5�f9�4��L�ҹ��sxm.t�ׯ�㤩�O;�3�M�Okpۦ����͍��ytb��7��9�G��Y7i�R�\#�4�� z5F�׈�YC]�A���JK5�o���������ڿA�@l�V��Ύx����8�u��01��;�T1��D�:�^?KQaZG��boE��sQ�[�*ž�ۀ�$&����(Z^ڸ�KY~b�����vd���E�JA�sUAL���b�U�?�X���1����ꑶ���%�[�{Z�B�r���bD��PM�:�pf5y�)u!?�<���(%%�����{n�PhN��:$�U�oy�ҥi��V���p��@P�������é�~bF�Q鹸�(7qT���o ��c�{���)���oo�g��(�X��2&�љy||<p�R?�ä�>orly6ǟ�m��KC�t��6�i?rZD@{44��Z���2�G�6��x��z9�{�	IqZŋ� ���mS#�v_��K��-�)���� My�ϐ�52zu��<r��,��)�*�����t9��x'�%�S��Þf�S�q/�>|K׉,6r�T�ԛ^#l�D��{a%�	��X( �bso�$4�<�v��ਸ਼>�k��Ƈy��W�fţ0��7��v�PeG��?u��"@s�pMe�$#���V��W��W�p�ib���@ӌA��<n�<蒙�<��un�R�?b`pp��c�`�~3�b[�ȍ�_5�B����lt
��Fx�s�����S��5q1��Gq0������.l���p�M�~����v�����v�h����H��)O��Ԥ��k�qd�8R��=���׷�999i�!q1��@+�0��0�OZyM������[B�W�>"���R���.����n���������̐��M�^��Xk[�_���}ɇMBnӞ��&a
<�)BHЪa L���"�Ef:222�*dTu|�a�d�m.�cb��O_����>7p��
���z���P\Gby�܏aH�����;g1�k]��sSF�n��[9^𻳍�E�������������N���[����TB��vd�K�x)ϸ���Wz�'c�R�t-�)�n*�"\�7_L��Ɍ���
W]�6-*�¬�@e���%�`��e�~�쫽,;l�|���A@�ؕ0���4��Vs;;!�'�C40��cȹ�ȭx3���]q_+kg/_�7�f8�X�ؼ��?��I�?4��A!��qUuw��u�#�@���Vh_P��)>��������Wc���O�b�7z�xo��vs�@��MS���0|m{c���~ܝ���?X�fSԽ'�V� ��Sb+�[l��oz}��a�F��7���'��w�o�),U�R�Vkp�^����L�kr:���Y5�l}�%A�w�2o)"(�mϣPק+Cp*
^���D�@AU~y���X�2ށ[ࣸM`f3l�(k=��%�F�HD���q�ϻ|�ڲ��R'H;S�D)٣�BC�NrE�bM7�8��#�x�� 8��y=0@��6k����㏂N��tAJGԏ����&�6(o!_��1Q0�'^���L	�j�'?Љ���e!�f��Ͷ-f|��ڝ��[�3سtW�����7��͍�q:���5ϰ�1�xb����|����޾�p!�]t�iѕ��,�  LQ2}[�n�� &��]^F�g�2G�	>?��x���m��
��M23|�����a��e�9�9 =z�63A�uY����wd<�����/v�cC�Gn�qU�'�ɖ��$��6��p��K�$+����;KBe��V�r<;��3o���������p����,˫
 o�"��0C�LU�?��I��X�gN9(Q|�(u��d`` ���h&,.,L���	I>�%^����}�OZ7�N��gl��	�7�?n�+@ N�\\��/��`����80����ϓb���Ǖ�YWa�/��һ�@��Ӝ��#�U1BZq��SI!
<�.�A���]]]ȧ�k��ѐ=�>�=�Lt^� }"�j�B�>M=c��1�H��9=9ɑ�rF�_�@���k��������E3�|w�ϻ�H�괙�M
�4;�}��w��?���W�5%��R���uww5e�X1���dN��NB�:N��ӧGI�H 9�1%A���-|��8*9x�D�r|PD�t2�v�G4���#�;�&NFg?�3)#
���66���:��\:$D<FX,�]�N����m�sI�{�]/�E /�*S-Dw�(�������aN��8;�����:��w(����P�6u6?�'��8���۱^��R窕?���3J�*���iA�E�&5��l�=\M�j��Q�"S�H.���D+�=#���L���,� ��쏁ϓ5��`[��7���=��r�:��� A�S���}��}�����p�x��)?�>y\di�ꋟ�G3�)v��H}O��C	�(.�gmvJ˝�i����ƟNk=��T\����#؇��ૠϊ���,�RC,��ZĴ� �����輸���X}�y@��<�<�Ҷ�;t�U�_� ֮Vr�.�p`�<���;%}���ggn,�4��������4/T\ry����w�}���lD2�d�щ���^���BG�k�t��驫�k�jjkC�����F��\
O��������%��Լ7���1q�k#�w'Jy	�rU*��ӡU$���d�X>������@�b�� ˵;��+���}Qc 0�U���]bB��<�{b
�cߩ��\�z��g�s�Yv~
|��o�xY�jOE��{݂��i6���_*����37z�D����+ A*cpu��m�P���Z{�m7DNؙR���e�A����hS���]�G�31�.a�1Y|�c�bcz~� �����A�k���Ϗ^9���Ҍp `w[�my4߽�V�6p��@x�4��;��L:?��.��8wg᪡���%ߴ�n�F�v6!��I�%/��t�B�����;�Sl�7�ѳ�R��:|���M��	��ޮ�u,��AI䵅�G7A#p�@��u�*FdeeY�|�w57ۉ�D9��&sV���7g"ڼ����dN����l<^uB�"9�788Q�YC�;�7�c��C�28)r����$7F�[��%�a�쥘+�`)U��8�o#��&�0��>~4� �ʓ4�'��$ܠ ����{��N_$�R�w|�u�`<#��5�y>I�\�!��|�~])��
���[��ꥄ�P�.~�{��_m팶�*C����y���[�;��x+�[+�OE��)�m���^���Tܗ�r�?���� �F��;yaN��Yˇ��@M��<^2�2�2얕�V2�?��T',f@K�;�,�}X\|�����ڄ�;����/�=>����Z=��D؏����u��	
Pj�k�"|;�aVdP���oMz����dN�,�_E�����ʻ��$Я��D�\Qt�̿(!?��}"�$�h�6��f.p"S�R�%�}�')���� ��8��D��"��}�2ۤC?�$B4Jt`�EC�5�a�9QFP���<��Dq�-m�*��Mz����#�vA+�*ȁ���ByŤ(v��o,��*��7H�z0.��nƷ	ߥ�o1�\�E��9��ӟN�RTr�Bo��9��cR��
�}��ϲr����z:Ν{�9l����h�}��bnzό�,1}sW���3]�'�óqGX������`蟒:�� ���app	�?h�p����0c�6ڗ��ၒ�>��q��a�	�i�V����˛���ˏ�~*��[�����6緟��11'nhc')�+Su(www�=���uS��e��ߛ����k������b����_��Ạ��
7e �o�����'͡�0�j�?rr�\N���x��Q���H�o�MJ5,,a�3����0[`���4�`γ�76��;Xdd����}�Qw�̠H�Mb��/�����?�=!UѨ���2Gh��aG(��w�Ve_��A���8�B$�]�J_@���tM��^X�e��͒�3�OP=����A�\��K�{����ӳה�6��q賞��oA>��q�&���yW,��B����!'�T{����B�
���o4��2�U�9[~[ҙ�a���ڲ�W�j�C��^��,_�4���b�^Xv�q*qD��[� �e���r|�G@��X��=?Y�SQ�ٲ��&� @�ѕe?��U�#�w�JA?�Z�D-ea5)�2���f��Ss%z�I�9���V:V��:%!»`j�]�A������ڧ�f[��k��&�q�e^�8sP��n����+��hi�O�c���Ǥh�F�Tz@���"Csa��j������9�ڐ��e� ��sA-���=�w�K�(����lAB�=�6�
���/d"�n����g���Iѽ�*�pE����L�����T�4C��Yz��GM%#���:c�v=�1�����}����q��|9�Դ��`Mc5���u�c`���)A��=kma�m��D���pX�N�گ�`�l�%��PK�t��=�����o���-"��a8�)j�	2��(��?|�ba�:�F� q6��K2�W͜�h����_�&wYx��9�^hg��a?��||zz�;����#�J����C5(Yd�h��"��f�����}�!�SN�@Oz�υ0�9�2r�_�"��#�a��v� 쳁�2����rV%Y�BS��s&uJX���~�?���u��������C��tx�1@a����(�0ʧ��U�_�x#"��K�Ǐ�qڀ����q��/����&����
��4�q��2(j�uI��ʈ�FK��_�3�D����L���p1ԭ�X�}�t��A(�YNR�����h���B��7ٚ�2��|�L�`^��#��H�}�;͊,eqLc�bΜ� �@z���m�:�\�&������7n}1,X�iS�73;���`6�777����yЈI�(��A�P'��z` Bҹ�9�h���&!F��B�X|Q �F҆#���u��BAA ��) �1�<.e2]jV�����V1�̎��
����=O��SMr�4=���L4B��V�%"�"�J��j� ��(�$�@UY#�^�
 bv�v-�-�����f!QV�/DQc��>�g���"��5��M�MӴmP��iCh��'A�IXĚG[���DNDĊ�u�o2* T��:S���`����|���,���@�r��%�.�p3�,�aˬ�����effP�D�.��ɉxRn�yb��U 22��'Dd*Z��7�{EQp�"� v��
��fq��OQ� �Q�":$�D��8&mC /= X�̠F��smh��Y;�p4�}�N�6���>@��{o��#:�Je�������9&��lL2���~�(+ IɄ��}]�����}F�{��, ,l�#)��o�-qqE�YT
*�����f����J�t%�)�ߑ?Ɯ�Prw7M�;el
ǊTO�h����`5�Y{c?D�n)z/nrqN���W����|<�8v2�������aU�eQ���5>e�»��ʲ���� �n	-n �q�����n??镜X��,��@�g8�-�}����{扢�0�%dG?�>O��F�&�m�9��D������P�c�5"X���QۛY #�#V��=��b�W�� �sD�G���W�,l��5$���`@��WC�<F�GcD�G��%D�!)����^>���y�=!?8jB3�4�/v�o�JQ:�~���k�JW�s!���_�|����77777��;����j�o&u#oQ�jV0H@��&��;m\�4H�� :���-n6'�&�إ݄@)|�Jp��c�?�:� �sh��=�ٲ��#jo���hK; �G}�
p�4��{J�S������H�����Ho,i{c҆`Q��{�����'MO�Y�����,`����b��#��*��m]�fEｋ�>DV6.��*���a"b��t��MO��9�拊96�vg<g"
`	��h]v"ɓ���E�%""��H⪴�բ�It|�s	�w�(����I���� ����sc��c�l�彈�{{{>X\Z\.z_����0��i�:�;�*�#�ު+,�@R������bo�@9�x����ť��B�47���y�TՒ.����-�4���f �]|�۞`�!�RQ6�/���K�
"9������#�m <��&�����Y��
�t��`�P�ŵr�y?:�e���gq�zeݟ�z/����	��H@����؜ń�
�Q�:������l~�5���Y��j�5A?	�G˟��^{��h4��z0���k1�1uoR"*��9?���4�q���@@��zt�}@��?�l��#z�gN�:}��9�пY��,ƒ���zg[<��MZ) **&&v�a�@1�i,~v5~�E��97�G$���;:���
��A	����_���Q�"�2�`� Y��Ȟ��N��z&�{j�i�Gm�v6��u�4m�4@ M��,5֪BD`[���(˧�/�?x�`4:������S{� ��� ,��dP���J��B�
�R�L�]���o�3���\��9Dj��d�IԡU��L�%��/��X�Z�d�\6�D���i��;2�'a �l1��6@v�Dմ�I�x̾���g
	s̺�
!����d|�0��UXGJD�%�yɅ@
 ̀�=�HӴ�90���H鋲*E�����-�}ᑀU��D@#��������D�;]��PU��D�A#e��s �	8��C1�t\a�H �}-���z篾dt�\�5I���n�c���6G�}Iڢ�:���������_x�����������0�����57����3B�Dd��5,!�<)�,R2SUYL�n�����7�S?kAĂ�&�?��RJ�ȼ�ObE�>���W���u�:*x�螬'�+���s`�l�W�EI�N�wv�!�q�t� �)���a䪐�h��4��E����2�O����&>��z�շBM;k4��$i���� �1ˮsP;E�Dv���[\�h���#��d2�WWW����LBۈ%"Y����y/bYz��CUcT��E]�+ ܪ�X�C��;��`���R�����s���R��i��}e��*����JI&)Lѫ��yJ�j���WUH�֓3;([:Z|=�3��yS h���\f��x�D�`��so>bǧsj�K�#Ve���b� �l�E<�r�\f��s�a���Z~c�����V��}j-U�Fξ��<����??�Nwvv�z�B�ݎ���:M�UU�jS7QE����ǴR�1�-θ�-�������&�� ��;`h,}ȣɑ,��/���G$I����C,
�Kc�=9
!ض ����[3��*+��i�~��`UM�q�..,���I������z)M������!��m��9A�j��
�b�=IX��,-��R�
1EFE}A�; �UXA�e (}!�b;�{�F_$��Π��%�Y�y�=Tr^N�j���sJ��q�:fE!BEdH�	�$:���{��6��r"�I�Rϙ������R��+�D�E�Va�$7A�,����Φ׮}v�ʕ7���S�<���;�}�����lgy9sw �;�{����:��W��m�X�۶�D �YBό��m���z~��������CD�̀�hT0\ƨZytT�;*X �T<�.A�o� ���~/l������q8�ݏW_p�0 `
��7�7NV��>y���%�t�N�D a�J�lןx[R"��c:�HۊF����v���0WYw��z�ˤ�(����2j1��^����������4u������X�eUU1M('�eYz�ںnR���D��BU8�P�H�A'�d:9��8��5��	��SZ��'x06��lɂ��X4�?C��u�$�x�^�q��v;">��]�sn;u�3�����s������e�?nn������i1�"'�EP` 4h+��9.ܻl�cg,�_#� "��C�
FR�?i�h,�F��n��
�́�l6cn�x����s��{VO�����%�`Aff�.ll\�=<<�q��t:����y��Zb>���������H�Z�@F��0�&i�!�MU��;��<��1���@Ĭ��f��9�*b�Ġj���yP���t�<�}"���`�ӊ|���h�\X�n��>>�>�����l#�K�;I
��"+���tKBEB���/.}Y�0(:׊� ly�
b(��J)��ST�s]G?�,}ͿOj��Btz�"��D|�dt���4rKt"�֎Y,�wC�a�w6Z,D��Hg������8s?����¹�a�R+5}]K���D*
U��o��F��t63�,�,�٬�~q���wc�f�A�����j��E�	8'�Y���� !�M����G���79��+@A��f-���)����G�KUu�a�x�e�9��A���sմ�ń��3�?مPU�scl90�Ke�=����h�
.ٚ���'��,�~j�J Ĭ�VK	0��!3s`�������G*s�%[>p'L���Tz03��������?al�Ln��h�sB��H_2u��v�:uq�8%K#��Ʃ�T���
�^[�<L{hAE�s�ɤm��p�ݧ�2sQT�ýmCh[�V� �#���1�S�A�-X"�����P���ԑ��}�tF���mۄG��=� ��+�����X�G=
E�t��
��Dt��Sl����}1YY���@�!h�͛���C�X�;����u���?�I_'�>vղ �|�?�Б"�&�#�@��ܞ_x?����_l=�r�-!��@��!�!D�%S��nݺs��l6��)v�X�U R� ��h7�z�% drNN�����i����c�����SrI�<`�q��P� Y�Ţ��D0��n� ȡ2�Sf˭�l7'*�Ӷ�_V��  &UP��H��ə9����I���i���Q��)��쬅tK��~4ˢe)�N�r���w�d����*?(K 	�^��9�Y�&ů����8�@�c.%�xH��,���|�溌�|�Rڹ��a"Q0���ɅS�qlB�.�,f[��,��?y�������|c�0���9�{+�w�O��p)� �H��!*F��������
�eQ��\�v��a����XeYmۊr۶��A�h�`�a��m[D2�!$%DH�K�'���6ܜl"��tz�ƍ�`8犲��I	�&�b�Js8б��y��4�����C9��O;�����#��X�c��HГ�}�z�`k#�,,A:����FU|������Ի�H�w\��'t��z|��U&)3 :R���;ؓ~��|�	}�=,c��%��Dz��'���I�̿Xo�
1�D�j� �KI�1���{��l��H���l:�V�W'��nۦn۠�9#=h����M�Y.�ז_�J���#�sˡ5�Y'��`�����~�)=����ﮓ�g_5Utb�:t���'t�ᱣ�����)v��vH��Z�|-k�=��\�T�~$"�s52D��t�]RLO�+ŝ��8��A刼�f�:��V<wM !"z��~������(9���CӶ�"$
*
��!�M�b"��}v���6�\U�V� 
��� M����Y"\<��\I��ݬ=�
T� ��CDT�:����ܵjM(E�+RK�WP��Y � r�=Z`��k��>�^M�*�+�K�ۡǶZ��1Ȕ�\�T����l��ˑA�7�a�iL ? �l.��EA�D�@�S�2 RY���4�{�j���#a�}�V�۪Y��U�G�H��t��1��y�������<�*�]�Dmܦ+��ر�2X5�,���R1���L�觰P�g�z�H>_���\��;��F �m��9FM��s#1��fEA���i{9 `��=���вs��;�EȊ�1VmA$�6��65�GG.�)13��mdɂ{#a�*g���<JU�;� �H4=�(�&G�eU�O��z	�'����)wBt�y�3m���|�bV�]hy�]�W�ݐ���X���eʷ�q�=W�{�(�#�KN$�6gߙT%"��J6%��_���X3N\ETB��y'4y�%�!i�
�.k�	nb�!��2�E��.�B�TO���]h� `��zƬ�/��T����4�\{�F���.�r0\h[17MS�eY���m�b�F�+y��SUB�	����s�U ����{�<�:򁃈�+h���E��q!�w����w�N����6��ĨN2�cv���đ�Z�v���]��� RcR3���w��Typݑ=E:���jz����`.�0|$"v'�Yv6@D?5q�hJƝ;��[�u��B|��2�b�;z_��Zڢ��lf�<0s @Ωj�4j��d�(f�SU�~ .=U�顪�Ɂ�P8� ��$"XQM=�57']d8ʻ%�C��l�-�n�QW5� ���ӳ���,g�HL��6XMH�sNTDY���U(���E%�S����4���E�z���9%b�]����u�b�ih�$��J�_�^[̕��q�0u~Ok�L�cA�b2Flrј�D=��o���-P�d���["Ҷ��`h����$��е y"g5�!� E6ǠFL!����|�$&,�ӔG�}APJ��nG{9Z��8�\X��&���$Tw�l-�r��%�2ᖥ���lV��A�!p��V���Q۶��m Qe6F45G4�%q���[_��m@	C��LT�g,F�"�����u3��D�*+ K�bU�D�E�`���i�<;Y �fRЅ��jrM��ۼ9獛�(
rX�{��S����uH�vS';֋Co�Zc����N����M=�p`��ڇϏ)-#9Ot+�"���"�#7�$��4f���zҸ����O�+��&>��<r3�bD�8����q�e7L�?/���ɩ6�ƺw��h):O�� D�`����j�e��8�6����|��"O��QEIS�q��@}1���v��/��9�s����JU�YBH�u�Y���O'	�f�4�h���I1.�[���{� ж-�N8�;�Y/���NUڶ)��c��I�|r�B(�j�9΃OӒ���~�#�}"�~ny#״*�r%��L��6��+E�3�n{;Ţ mk�~
}D����'����m4���D��|^�OF�&�S�����6�~���q#�����# �"�B�9;'�U2�A/
�)A�,KQ��1,��K�������ChBh�G�޶M��ꈒ�FU%	��T�1�&L�>M���H
Q䄂�)��*����@v�a�AH��$�y���2� ���J�	)]��N�,�<��DDu]u/�ڶ!������@�#���!X����B�lE��ass�!։b�S���<9O��}�϶nِԆ�AJ�4�"���V�h0,Y�@Tf�W��[k��aQ�HԔ�� $4�X�8�l�e�2e�v�c��sVL�*�"
H&�֓)TJ.����]�yw3�G7e�sz�����:h[5����X�<�P�E`U�Ȯ-���U�֑�x:�8rUYB[7����h�S��ޢm۶UY��֐@,�ZX)n�5J��z����TX�< �J1�d��ʲt�~IdS���h�`�L@�舢qc�S�j����}�� BX�5����y:�����F� 6��t�[u[v�����f���l���&��4M�)W�3{��{ADR��d9����lg��}�#W�젪]6�	`G7��1�wF>�LlR	tOł�>\�J&�5Q�Em�=rF��E��}^nX�bTP�M[%�B,]��(�a�9�d_D8�u������l]m������1�l6���6�6G��4��s+t�+�Fܘ�jdx����U~,/-��d2	���(P0��(���MgEY�uc�a�-W0������~�e�����n��9������uvVk`��O���0���(���:e���y�����b�w�8����z��H�c��+��fzY��@��I���K]���ٵ�=P�� "T	�F �^9@H�gQBL0#���
(]V���;�!i�������&�TDB`f�ݒsa�X��C @��F�NS��[��q�:��K�^�Tb�F`�D�g=���o]w��3 �_�"Hh%$��$�!Af�F����1↉���B-�������N�����C�  �"*�З�w��7V�C�l� ��6��sޣ���g!�j��
3�#Rfq�D8��6� ��t�&?����c[�Z8u~��H:C8�g�<E���FciO���dHGZ���D�6Ĝf���H*�4��E�=1��YT�m[U��!��-�9uh���T3�!6N4K�ޫBZk�B@�L\���W�Z$��`�,KKC_z+95���a4� ��d�I[AQ��jQ&(��Dr�'rEQX^"v�-K3��f�b˶T�� 0�粳����o������j�۲�H_JY�)�#�E��2r�q�y��.Z5���e�Y*��$��ʘ+��4��S�#�_��m�;�������d�%�pB��Q �I.4�9����i���Ėm䀺�ˉ���, 羙8��u��}WS!A�����8��������&� aQ����{���r�/�������eYF|K@��mCeTꞕ���)��#r �&�-�c����1>pKD���k_{�{wppp��������G��m������҅��++Α�����񃭭�.�6�)/�����Sͨӏwgj��?� �������������^�%�X!��Uea ��H0�E$r1$�f�V��j�.̐_	���{Ѯ֬{�n>"Rha��~�޳����s$ҩ�޼v^�e�QF$�H�ѻ������$8cYt&R]�Õ"�\�x�s��h2ׅĚ���(
@ �1����ȱh�͔US8�(�⒩�I%����h����TQ���Hj�T�ME�0c�7t��`�n)����A��8J��#�	{� �>�>D��v{�ݍ5��6�q��ݜ�5�d1� �L�mA��H�10���	X[kD$QD��Ѹm1��T5�q�-rm�Q��<	ز��QUrH���G�E���:�ӄN��ʪ�I"r@)�R��m&� ��� @y2*����!�-�C��l���-�P C�"���EؠiD,�2�`r�0��n��`vD��h.Ԡ�X�i�V���j�8�1怨�`�)�!��tZ���G�+��T,��'&l���j�5����z�S9��~�G���"!�@._5v!��9���U5���{��Oܚ[�qL�U &���G.�1ĸ��*�o�`��,U �q	9e	MS�s�X؋�.V�[��e�&���:4�7L!e��^g�u;-{�Q&�o�a&�8�mX�d��?��س=j^��L@@G'쐾ȶ�L�s�3�B��=Ի�M!�Lb��ι������]]����Bk�Y��
F  63A�Y�EU��Tr��t{��$ǒ��s
�"�tv���_ܸ��o���ݽ���#D!�/��i����?�㧞z���vዋ/^�~������,MUi�c�v���h�~�E���J��X�C�4@Īڹ`eB G�����h��1DCh��9�&���IuW	"ҹ9���1[&;��Li��	9�C H\A`Pk�*cC��K��C��&�M>���xt��h��^e"͏Y	�s_���)��*.%��
ڥ�y����نHM1�%��s���tmԼ�MsR�D��]kŇ�2k��`y��̱#.@-�b̒E:�D�U�;�D<��d�$"�Ɓ� E80�E��CQaV�M��vޙ��B�����su=��P�!������V%*�K��I=Mn��aǴ702�:K����4���C���0T�$!�Zn���M�e5l��iZE��T�9���*BhC(���#�#{��Q��t��e/���j!#F��D�6����	N��@jC
��R������k�4a�}x�6���>��{ r�-�+���ߖt������pcc�{?����paqaqa�����l�E9�`���K;�LT�ж �'�0�����w��#e����m�s��*�B�]�J���J,�h�}�Y���T�i�F��8F�I���}����ދ���0s���x�Vl����K�AMI�ɲ�'5��#�ϸKY٩[;�V�dZ����={�9���y������O�ӭ���m		9r&ɑ�ڶ�ճ��E���2p���Y�&z��b z�ͺ�;��"�"Z}e�7�},iP�r�l?pw�;�$�z����54�����}���A� X���ʰ&��=���R9q3:<'m"��n��Y�=4m�Dm�Z�b
��a�>�Yz;`r�i����r�r�_��ha9@�8���������������ˋK��m[U�I�V�G�F�//����9����loo�Fc����Sd�0�F��b91҇��f:r�{���ӗ �'8��?��k������WVW� ��3gϭ���t:�P?z�p�0x��gU��ϯ߿/�BD����"� j@ ��69`�_��	ީpr���f��87-I���S��;(�c���
�`!8��.�����9� ���$BU�d-�� �ZOH�AX8�@����]_�{D��;QenE��>��lrRm� �Kf�3�ζ%�"�j
Q 2�%�9�<�5�e�I�*�0�l3w��mp��TU�9 :��~6�C\ᄨ�^�p�nDE%������ii6�"R���f�^���UDfh���$��B׈	?������1����`�z����F�FR"l
�,���\[�Eᓍ ��Z4�Rp�c)�/}�o�&��;z�	I;�FE�9���m�[U�:)���As����̀��Qg�M����M�hస���E��),30!ǩ�RƘɿk3 �ݶ�"#�Xۜ���ՠj�&� ���_{��Ñ�����d2��ݝN��������Ѭ>I�����i��pHD��(^]Y��Kn`��D��ta��G�9H��XF��$m ,Q�XTH;��,Ԟ����_�dEFB�R���sBd���qE�ⷹ��
��.��T���W�4E��2�˲���İX�� ����L�GNI�sW�^]^^��z�����������/_>����y_����gM�  �h�ۢ(���U���ظpFD&�qhۦ�e��v��ƓqbQ���R*�>���R9�5E����S~)���7�.9U]��!R<�*���'��f ::��Y�B���PN_E[��=�{t�{hƘT�r���RwQUU�rppp�ܹ�,��G��h5xD�0�d7DGC�O}��"��r�m+9W �!�Dd��)-Ｊ�677���/\�P��[������,�BĪ����_���X��W�.~�˟��{xx��þD�s>:ƽ���9(ho����IXUR^'å7M�ރcE�T!B��1Mc���9��:SQk�ܶ����^x����Օ���������������Kˋgή^ܸ�Tdoow_D� �(K��+TXʢX__w΍ƣ�(�����~aq8�NǓ�ʜi����]\�?\U�=P(M�f�	ck ��a�i�U�T��F��� Ή ��y��VVs�X�ŋ�hԐ�@����p�6����#��ͭ���x�"Q�@��U�C�IwD ���3m]L,�F��Ǵ�,��Y�?Z�
��KKK�MӮ��\8�.�8��|�������K�����������3&�����E�4n1�t�;�,��� ;���;�Zn�氥�Em�ڝ�ޅm��̀�ȚqO,����`vǧ3l� AMi�X��"�/C�S�U56�UU�=��QG9"h-�DD��8eD(zD�b~@(�!p���d%�y��>�O���G�"RFH�,ʮpH@�*M��j�!�e%槙%j�fUB�`���w���1��DZZZ�|�������+_�����`0*J���|���4������@���z�����ٳg9�ݻwg��r��p0|���Z&b���^�B�"�� R�P�.�G)�h�1d���G^��t䐐�U� M�+ƄiLa�yf
 `E�v`N��S�$U!�y�lM[���,�-�5�`�E@���
lcM?aT hQl % ������$���6����҅�����3gά��f �z����҃[��@D�s� �f������i��W��՗_~i4����/�������W�����C;=�5��*��7�$ *���2D��Ot�6 ������&XM8`��?�!�,�h��Az���F��^�m�6&�s&i�
��%-9�s#��i/��;s��ֈ �����t�
�y"����­�0��\�)��8���*B�l���Hۆ�,T}��W�"�'@u��"r��f^^^"�=|x��m��W�� ��Ν[���/���9���ɏ�_��,+@�)4�[#��H�^���Ȼ'I�M�bN��tLO�!D�/��c|6���7	AK
Q�/]&��(˅�P��)K���ZU��mV�WVΞ)��AAˢU#@G��y��7^�m۽���Օ���w�ί=z�����ooo���9Q��q4'ߒգ��c� �3}���#�Gdq��җ.A�Y�n2BB�:ǲ7�V����I0+Fh*"�@I�!F�� L�!�J�c��`$�1��R�Qk�( ��O2�B�ۈ�KcBrѬĔz�RC���%�;�5�!��!����76.��l_�r��w���l<>Dt��~-����o?��3?��_��<�TBQq�l�����j00�n6���`9(L�O�c)\|�>��U�{����^�mE����Iƶ2�E���d�_��z��{�Mo����L����QBh��RR����	�.�jʍR�"ZD�-�����j��+ ��Ҷ�'WU���E�!K�׾S�2Z��CI����	������.I�(m�l��Y�Z����|�����YB��MH�,���i����i�8k}}}:��B�Y=�LU���t�޽ݝ=�O��h��A�0���;{���G�/_��>!^�t���{����l�MC��;'"��tqq�n[��svK�K6��Վ<�X
A��h�ń�ct�yB�s�Ԁ�L	
2��#��t𧡪#�	��o����e����^�G�B32��<�s�8D��[��~�� �r06�Hnj���Rp8�h2z�왗^z��F�â��{_�����|���nݺeI��X��#K��F�����~��&��}�9t�|��+�}�������{��=|�(.� �w����v�K1tT`a���"�J� 	�=yf�ĉA�S�LQL�GH7O�n'U/������V���s�N�W�7f��f�z6+�TC˖j����D�wZ�3� T��D�}RPA����m��M]������t6��ʢX\\��mhYxye	 ����fv��?��������E��*C� ᓏ?^��;�aYU�?SU�ݳ�����	 ۦEG��y:"��l�}FÓ""�Aʧh��݌�s�|�F8�G�d�FČ�����������t���]~2M�# m�f4?��TV�t6k�6Y�ѯPU_�m��9s�W^^Y]�}��t6[\Z|�����G�VW�������7�u��%B@�T�t��ݞS�c�9Q>�o�y@U����O����sH$��E�rB�<�ʣ��_#::&LT������$o���Q�1Q;�w�jڶea�gv���"�M�\�Ή���֒�3�����VVVB൵s���j���2\��_�t��gϮ��)�EG� ^�l�	���������z����۷�z�)Um��է����w߽��E 2�0���w�CpK˪ �!�i���3ƺ�IH�ѱ�,ϺD�W?#��@�4���(��B"�\׵%���=f!r�����,�2�LD�+%٪M�s�s�,K��2\LA��QP�g��)W��K{�ҷH�M����*��
�"�e�Z(���1
���3]EDK�V��{���UA�.A���í��g�}�����?����J۶;;�++����(��i��,�V�.���"�h&�=���ٵ~�[�o��ʫ��G�hk���я��)������{_�%""�s.�at3Y�%�&ܥ�抙8ҟ�^�u�5#�%�&2��_m��9$�� 
�& �Y`�ڨ'g��6F ��om!牾�e+n۠��$�ӑ���z�,�t�rA����T��)�E���<x�pg{�ѣ�����4MQ��zF�.����w��M�Q*�ƆV@Ӥ��"r����?�|qi����`P-..�+au8\`f$�'d��K˜_d�@r]Q! �I�:������_���	I�q<�����0�e�1J�75_n�Y�&�Z��_������.�Cl� jT���j�v�\�67T$���}$��0�_z����������_��_]8����v��ݿ��U�O������j2����?{�̟��_l�l���[W�\��~|��篾����~�W���o���W��~��>��Ov�ҥ��ַF�ѽ�w<zԽ"�"�(�����`���?�LVVV��j�z4�L�S�Ø�/�+"�p0$G�b"�-@O.|م)�����*���u��_6�"��s��h�ڧ�^�ti:�ܾ}����'�I]7�+�ۻ;��>|x��ϧ�I?l�v�pEQTU5�677,'dyyyk������j@����}��Tʦ89`=gnb�����1ir�,��VT���G��_����E �'�؝�_2��Ͱ�`M��6��_���KW����[��VU�K�P�ğ���@L�J�v
�1�nJ&��)�s�id�!$�~b��&#5��,R�)��́���S�Dd<� �իWVVV̯��f6�y�s�[[��o?z�����5mCH96m��&:��|�+O=���[���G�����w��������ynkkk<	rY��{��K�`f��"�w�$^,E 0v�\�3'���Y\D��i��8��|i�	`���,��H��9m��m[f13�R��0�<�* ��`@��h�B��*f	ªZ���X��9aaD,�JUY�9�ĭ�B��,��+=���s�B�d��q����f68GH(��G9nL��6�#�>��Kum� (�)ht�ƍ��݇���E�k��{WU�lV;��l6���{k�#!�,�LKy皶������t2]]]�L&���x��͛7��,Kq�"(��d2!2��s�:D�E�ͥ)�0E�7�G�
873��ʔL�����*��JF ���^'��+ʲLR��hj�/��_*�����I�v�(VL���$�%�Hk����\�9�Ű���NZV�`0h�����o߾=����Ȼ奥��6M���� �l�}�țm�#���*�������������n[��L33w������D&A�,U��&Uu�z�^ZKKZ���Z?Bk���b�"Y$H� 	d"'d��;�y��nfz0�ر�=73�"�
����!�s��>�,�6�n>�j�͓��?ݿ�Z\\��i�C|�c��}0k;(���;����a���K���z��5�2�Ɲ5�v3��$˝χ�c��S��L��N�[�U���'�({�tl�J^3FDĉ�jb;,^/���}õ���X!s���٩��_����������Φ���P�����?z��������˽�����6�����{�������ɳ��������^<�����������ڟ����߿�?�O��������O�������c�������K-p��fս��������}7��������}���qғ�'���׋��R� ��SL��3�w�bv�l�<I8X"F��O�~`E$�l���UI��z`Ŭ�E�i����)�����g�*�W��z�^�c����AT�EJ�i���{o6b�:�����_}��7�޽7�L./���/�b�^UU�����g��`�fᖭa	�m>_��ψ�{��TNy��~���
�����;�(}c7Ashw��W.4A�q�f*�
1:�z�r1&s�#f�jZ�f_ K A���QU�i����"
�sC3�a7�3FK��׆��Y]<{�*����''/_����[o=}���%V��f��G��b�X|�٧�������Rv�KQU��tq~���7M���7��JE��E����~ҴM�*D��)�X��6�Z������H��rRZy�8q��y�^�  ��ȕ�F*@-��O� !�\,͂�v�@N:��0[�������S�y�I���#�#�W�ÃC�^���������z�ɏ��Kr˵�<˝�$�Se���٭��,��c��Y1N{y��V�zs��ک|�`�+*Ѷt�����i�^GNu]IJ�,�xvvf���Mӄ���mۤ��zd<��zm���ZkB	7-������ج�����?���_�ѭc.U��F��l���FW���\��PB�(�f^sep�H兲Ev��g�]���Gf����Ǎn��Ck�0�l�|3;��=Rin6��rQb���Q/�<��ˁ��[ �U������5�XX�w����c�1�.v*Z��ꨮ�k���M�""�7��d������Զ�z�j6��y9�
Z�DE��gϞ������{�>�����~<�����/>��_�2(P����2�ՊZa�����yaٳ8p��5<|s�� [gb�i�l���~�Z����R�����:w��\���_�dTC?�N�T��꺮�kQUm�ӎ�=Њ�ގ�$�W(9R8;?{��Q��7�˫��r�u-������(s���X���c{~q�Z.������'��y�n��N�>����k۫��'_���;OޓH"5�0��x�����qLq6ۻ{�^�����{o�P��F�i�v޻�t:
>Ĕ�޹svv�ӟ��|1'k�1h����y; �wɇ��Oz����S�!�Mw�l�)&�!u]GH��%�i���ͦ#�s�ͦm���d��q�9���l6���[o��_�׿���mo�:�w����u\�_�R��%��"0@��4�����!!]����!]CDr2�0�z�{��ٿ{v�}_��}��sW�XwE�닗�����K�q������ub��5�5���x��G2�6��B�����"=�.�,ڧ�9�d].uWh�i��M@`�I=�آ{=y����5������߃��D�����|Lʄ2H����2ߝ0�b^��w�53�OF���������؆_���!�w��rN_���湽AS�o�2i-�|��;�Աݍ��w�k��m8���Ov)XDX��,����i���~.��Џ�� ��X����<�	-��n{k��^�U*��C]�@m+ix���T���	Z�(����÷�l��z�~����O�˖��;��g�S�h)4��z��Ә�d��7+aᴴt�.��� �� ����i��FR	�zǆ�^j�K���4�HP�°X��C��mۡ��$M�%��K���]��}r�l��CB�5��n&<�/��c�{U��d���f31>�t��߯�f���3I���TMq���Mz���)��#��^�w7ªN�j��2�O����{�#�m�(� ��gJ��B�;<7�f%��^�0�I��d��z����N��_����;4��\��,Fs�"�쏄W4yؒ�����?���h��(���'s�W���} �z�{"LDou���ػ�Hl�|�3��j.�����>uEU$S�m��3~0��k�6��\�񡰗�U���%!�v_,u��Ye~s�J/�=Z�$V��DBI:�p+H����O�4�A/��]n;����q���c����  w�{��{e���?-�- �Wf ����cc�al�.��8n���1��C���:v��r�c)3E�ཟ�A؏�&h�{�d��q��ߝ��
7Yu]a4L�W'�w�M��(�]5�}���dA��^��T��������賬R���q�����#�{}��3���Q��HiIqq���Ȉ�͌u���ؘ&[D�HG����[�,9[Iqi],��c��8@wD^ikt�G��wK���*�[�g:��EZ��G!�s��GΥ�AQ�b����l^.�_���7D����|OUq�(=_-��pE�=e�]�U�|�����A���Ҝ���ҔG�3��\x.0R�iZb�B�}B/��9��BÙ����m��塦����������ꅁ����b
{�N5��R�]hp��r�d�Xmz�X���?���j���`M����Y�@�C��Ne�%�T�#@�0&�2dߔU+����y������C3�sc�����f�Ay^����\��v�G���R�#��f%�,�";��@�V����ϐ@^�^�ղ`��o7��[�a��󵣿c�kG�,�ìΪ+��BH��q�������sˊ���_]S,�7-�_!o�����իƠKG�W`�d�f��֥�/Ε8�� 3�13++S�qE�Z��6��rؕ��.�|��`j�J �X��\324  M� �;?F�t$xw�4��U��	�^�ݠѶbC��A@�G�jH��PU�M�X�Y���e6�¼���Ae��KG
�ޗ��a��[�4&i:����b�I��wWw��7�J�R��M�x��&�{ �I����L�d��0������Э����� �#��L�r��[
wW�i��2ŷ�ql�/�~.9�FEE|3���W�w�F�������G�������p�p��VQ�O٭�U�9�A{�����ػ��3b��(Y���e�j��C������k�u�1�L�����UQ�(����2� ���­E���yP?F/w������w^�`�P�N&�A�ۛ?��q������8����ڰ8����:�ǲ]#�qtz�����A��##;v@kA:hR>v��b��ݍԟ�����6ׂ���������˩����������VE�ZR�<O�eJQ��L�:G�=}��OH�9T���j�;4��%LЪ��83�
pI���)Fs�F�(�y�6;�wVl~��7�;��,�(��a���7gp�E΀�@��c��҇,�ł�
|Zo��N���퓍Tô�{��f6vv�H�-������.'��y���o�~�騕��-d͸����B;-��b�8k���ӆ����d	CnFX%�[������G��B�*!��(�
'\$��}����S����"nIO�׀͐R���C�����4�GݞP9Ø{�R���/�����8\I!gF��?�V�;�)�Q��1�i�N\��}s~t�K����߽�=g�����I}��x��vp��՟�..z��(TGg�1z\#��uI�y�k�������ʨ\�'*Fm�;�d�����<��Q!�QN!�-~%�t���%��hg�ģ�D��u)c��\�ɗ���� ���\ ���6������y�E���)�&��6('?C�l�3��]��s�&\�T)K�I�����[��s{��~�~�bGڳ��@��������|�'����B�0o�U������tJ�d����'ժG6+WA��@�E[98�݂���L����NRQ2�-�����blF�p� �all|uu�n�������w)���iՠn�&�φ'���'V����U�_jژ�mD���x]ڸ0Իy��)P�T3�`~��U�g�R7�$*%�P�[�++�@O�i	�AĚ�ƩT�P����Q���{�O�E�����vo�±���8.����)�K��3�*h.��4{���'nP�w��0%��UC��ٕ�{���9lԽ�������|5<�����|�hA\v�@����{��[��Y�8����H@{KKpD�\�Pt4������@FYs�N���Z�l��� nn���!d 1^��@��E�z�H�ж͢��?h���K?����Gm���]:�ܣ�ƗL���D�EFƈy�Z�E'6���Ö/���OP(�?�+��	Ч/�n��	a]-o4�̋��	h�#2��C{��g�4�Jݏ�;P��碿��%F��_��.1�h^z�h���īVJ||�[�Y�j�`�c�ȸ������ӂ��MP�uwg�蹼����8�l��30E^�����qaoW��Su�!2��w�������)�����0e0�7����Q��K��
wT�+�JFw�����x#E�J_p����r>;߈��>J�[���:�r�^u��OK�@�1���ٖ_�e���:
��;�4=�ޟ՘J�u<0KPp�H�\6r����u8J���8��U�U���ѡ�f��@��O���؀
/�!I��&=B�E�0?�����ȭUJf���@�������2�O"'_��(Bw#[�/�S+z�� o�
�;n%*p�t��7I���{^���n��۳��Q�y�߾����́\����v633"��U�4�|W6<d
'�J������LD�i�إ�1����H���R�1�H��k�SS�=�E�G3�i����ߦ	�S	�EM��޾��� ���^~GHW�,-�m�6N�z㮠���������=;pQ{���-�����]La;)N)�f�P)t�	N�+++ѡ�O8�9�9�d���~�0�""l&\����c+�+��(˾�#�����t��6b���x�B�ԏ�O�/A?�}��g���*���q~↜���CX>����u���Tt����tJ�g�(�?������$Rf�=�(t�2�$�t-���p�m�.Ƨ�|�V6�������'6?�I^N�z�<����dk�s��]u2���0�������b�6$���@���`0�r���C�������E_�F�H��be޻[�#�{��'���W7�h�ќ��ɘ��)�F��@.����8S���Jo3O:�2AL�uf�Q��쫚?����
,���Wy��`H�*��{��䉋�ȸC��T�⡼a/I���r2��J��@S�³�ĝOJ�ͨ�<�?M4���z�s�(O`�����d\�|������
0w�?.LY�-�K�R� �/��(���(/+�� /���pV�LW��O�V�Y4ʲe�������QY{^������9*���)�}>�!^�wdeM���M�o��5))L[���Vqr���vK������VB '~��c���!�?2]�---h��4�ʾ���r�PV�̬Pa�eDTh(�p✜lʘ>�S"�
��8|���e�|�ݝ7���������=����Iޟ�!�GBs����G�������9�����>��wƻ��@e�t���{i������ם���}��Ԛ6��>Ctw+"��/l�Ո��+k!�� |n����t����F�@�]�=�+��C��NӁBό�&¹|�|�v���@��t�3���³����r�jE|��E�����Q���O[$1���z�֤5�Ϳҵ�r���:)"��Dz��z�8���U���5ݙ��nC�}O
�����ۅ��2uykCv��)[lnO��L����|�s�3{�>Yd
���s,���%;����������z�z2mA`~i�[��-�Q�r��f��C��^���"n��>���d�A(���?m�i��3��ZƄ���� �L;�Ti���>�)��U�|v�o}ǭ��ٙ���A/b-�e0�!����Jq"s]<.3��}v4d���}&	蒋��ؾ����Q�H����ߧ�����>��TpqRv���:ֻ,��2��ȕY�k8��̾D��o/88�C�S��50X��:���� 2����SMذZ�[��dQ���F��ؘ���o?\ӂ���� }�$�D4-033G*�FP|��Ve�zyyy�hZ��#:[]P�	��)�M��
[��j�j�bECy�=���b(`~�徱�f�}�|�sK"�Fi$������hx+�C�c� �X����7W3J�FP�~������o?Po�S����^�&�B'Ă����!^��l��#���@z����	Tz������^���H�=d^Z0�fo��l�������6��^A=�9�=��aZ�t꧜@]���՗�I��������+IΒ��?�ѓ������j1�""*�⬩|���j�D�Y����S��8��/���P��4����L�3dL�k'�J~.HU�L&P8�7���8�$TQ[���b��u��=��5%����n�Ɠ�N�PU��+���ˏ
4>�lթI^VVa^��m���dc����o�us�3�f����]��<�)�z����冭V�u���
��7��j��PF%ߦԶt�8%����Gu�l��y�|@`Z@F�;�o�e�W�5�x=�(�ɜ���-��Tx��b��IȒ�utJ��e�'��<̬�6�o飽<o�E����֐��+��~��K�	k��3)�5oę$;�#�B�z�/BG�+��c��l��Y:�p/��xz��v�/���.�Y��8뺩�����G61!C�������b�˻��( ��� �&/M�]eVU��/�(��� ��
��L8�~��s.mWF���)|ċ�Z��)� �������5��<*�W{yo����_ba8
N�NM-\��>J]���^���Yy]7���v��o�l��R`pjZz:�f<�s�k�8��0�F����W��椇8�j"W��`��e����o2�zZ�5�m��3h���W���$O�'��-�>*x�I�48��DR�O��L܎#ｧ8�l�%�.���-��+p�Yȉ��:ǡ�P}��>IF9���/�1#����t�;i�q�}�h�3hp�},/����:�PF���꺢p~6li�)����nC� tq~!�y���O���y��i�B�zl��Z�B`���Z5�i�p��b����J>�k�I�f��R�
�F*�(�x�gϪ>���&P|���۶護�5��]y��u
�?�W�c�����n9�t����ym�mi��c?�;��?p��t�_���e�3�9el���?�mUg��k�����OU-��]N�Mz�i�Y��Vl�d��9����v�Fܜ��F�`�7}0�< �H�s���=�t��4}(��̫	lQ�aue��<����QSy�mm��뼥�́˜���~L��p��;��<�g�3�ʅʱ��X��a*\�}��ŋ��\�/
�K��Q�NM�j`�7�J�/�1MJ���{�4s����Q/������:{o'f�C
bl�`!;��2)�����L@��* ��'n���zʔ�RnM�I���	�f�:�@K��,L&�p��.�m�T<�s��a.���M�3���QD�*f�h-�Q2T���c�i��ξ�o�ݘ2|�����M31E���*���ڡ���u��;q�g�����|��~3�%��I�&0� ���K���ټU�PJ�}l�:�u��J��[��+�����8��z��h5�����S�	�M����rN`cc�|"H�[B���߮.6O� D!q9�)�%c�7aA_K+��)<�v�`h�Io{��.�$��%�8�"g>0�H:ަx<#i����uK�}��v�G���0]_;����k\H�n��#� ����+�,��P�6���͓K��6�	"J5���y!/_�R��;y���h���fac�x7�p�Tz�G�}��o�F��	dM��]k	�$yq2y�mV�l��n��Z ��O��Y�K�����\1Z4��LO�o"��|���X����F��\Y�������Gʮ^ʒ]�L������	���I�������X����:r��E�!/(C/W�p;Ѧ�����%��w��l��עW�Y�����%�ӕ��Iz��t޵�}Tkw�:(!AMMm�+8yMٙ�Y��i�߿.�
aw7���jY���/�N�qI)���T����ۍ~ ��0n#��O�����	�����׽󥝖8��Ƚ�!�+R����ه~�PtJ��95ٮ辝����;F�b�&�N`*�ʨ@�4���[k1�4Vr��ӂ;���D��Kn���V�L��d�X�?~�x��l�d8}��ݾ��%	�*�ua<�pz'%?w�ÍXJk��y�p���ieS~���VQy]䚩�N�Μ^���4 KaR=#����j�d5#9�� �������uma� ot��>�w��gV:�`�oR���+������q\��X�������������T��� K$� ��"���q�q�yu||< ٪t�[F��C��[G�����s]�@Ά�������D�Uxx�e�u�_6�0��v��T�#!vX���0��j	j8��握��k��=|���Ty|#m���{�=\l���Zbѭ��p���q��p�u�i�����1ڻ�aʷ���� �\�cDa�&޾��2�A���+"9���K�EX���;�K
���cL���{������q�h�-��W;ƴ9!���ǆ��q���m�3���Zp`:�S䟶�s����c"X4���8�PYո qq�d^7�7��%g��߸���(A��wY,������=��������qRnҘ�eM�y�{��$�B4�<L�SAe,&�y�I�������e�bBk�����׉Z(Nsf�4�sry������u��Y�������+]<�{<����m�W�k���fWT�O�G�\A�g�Y]������>��O��sd��t;#!�3=�g�W-zdؚ�&�į�m��9��6n�N9�r��3c��0`yrϰiY�c�RW��:��O�QJBzE%C�KT�2����qS>4��+�R�*�:�E��	�K�mm����x�4Zi]�Pk�m"�u�����+�W�iךfffAW�f�}���8��YXCXI&`�"X6�`O���-�����>�M����^�� d?�u�}B+�����81
ȴ�B�ӫD���H��k!�s*����V����{��O��S5	���s(ȟ�K�jF�K��	�u8ef�ޟ�]p�18���a�G�gn��-$�)��'~[��k��i�&��,��
��=g��`Z�c�x
}����ӽ����"�*���6N	1G�⧪������Rf��w0h0��vL�W���wXV���.�̷�K����QӰ< ��.���w���x����`�ڿ�E�E;��D;s����Dر��^Y�까}�L#|��3;G��.l�\ĺ�53� S�I2�u4;u�=��ճ��j'w}2i�
����4�RXZ��m�٢�Aw_{�32�92�%���%x�	�������\�J��P�&D{-����x
�s��_$��n�j����1�v^��H�u%Uz���*~8��2jN�����7�T���Π-�)��$�ڬ¾��cl��V���B��H��1aDH�hW��,�p{���J��^���co9ֺ�1��ڹB���Fׂ�
K!c�A����Q'��ODD�Uݤ0�DNNF��[z��>�6���@�X�<�,wl�C�B`�>�|F|��W�;�]R7<�|�'"^f�xU���r|*�#��uii)�5�d�2{o�Y���>�qy}}M���l4s���e��t��4��I�,������M����_�[GP 1��JyZ��Wv/�H��$���>���U�}.��N�z-�JTD>��Z��?�@��~�_��M����OW�����E�y��w�G�E_[/2��ñڨ �����u���G�������T`ߔjO٧oJ��u�تr����\{qĠ��^p���y�����#�h���Ӆh��`@�]���ޓ�gْ�^6LHt�7�*�
�2S�
�aD���bO���Yi	Y9i9i�YL��	��#��~��"��ehy��g������)�L"����-	��m�9=�����X{0!%`�096Q��D��D��j�0���e3��sb�{�� a�ϩE�~�?�Z��>O.���C��,#��`h�U].�C��n���"�`M/&������,�h�씑���������[;;�/����Z�#�������*ܒ��۲�_x͛�_�π�Ã�ʚ�{�������^��q[�Zn/�pw����Ӣ����lk�o$(	�G��n�	��ڒz�IcMT�"5F�uJ���F���P�+�g���A��O�6w4�����*Ƨ�U�QfF��*�k*Z�U���M]y�vU��m  �gW&����L9���؛���������G6X�*D��"��g�88E.ɶ�b6�լ=Qp�Yc�SZ�\���m����W�.������}�1?�M�6���F�K��K��T�O�`ʉމ����-9��m�e�چ�ϋ�)}��~r�Sf\�"�J��]R�)(��fUr����h4td<�R��
�K�ݱ:��+"�-��)�_��<��qv�Sz3�E�H�Q�p� �}�qbM��=�i��jI�GQ,��&o�}l7[���s��*����f~�Q�V;��@�8�0cD$?�=��
:o���1�́\��᜻�=��$S�80�i��؇"�*L&`*��gP8�F�룆�.��d��#@��e���2G�v4j&L�z�Lj��L�N�n��\Z�;�,�j��'E���������ք��NN����2/���u�:s�����?e��`�+hi�ܷ�~;�[�oY_��2i!X��Sb��@�%��v�H@����<�^��b���J�`�}N���I6�>Ek��J�YyYpoG��Y黶Q+OZ���OI������2����Dy�@')��p��*Os�(l8�S�PG��g��4��+�����|`�D�k����&]��ԏ��Ke�m�;
�K*��qUbPx�%��t�7!�}k}q/�u~��fg^xI@��cx��S��٠��N���ylE�v�������&�˲��m�k�����P�Ĝ�&�k���*NZ�&�1rP��c>4ֵ%٧��4�yWd�_�ޱ��W2~5෿��:r?�I���g`-�{�S <bO�n�u�a�|�O?�՛���E�B��"�����Y�(�!��B_�);�-�C4��#���"��s���+�7yoU��'h�raB-�����ҝlԘYGm؉u�_ o�/��<7�;�;�:;+G�g�#�l�/���fv�4��B 'o��E�S�kʄ��-�w�B_Z4l��ĳ!���Y/�6W��v���7�"�5d/t��.��e��G�Bl&n�xA����o8?~�>L�l�H Z���[��f�90��>����,(F@�L��s$!(+�ң`V��L(W�����N������^`�S*���ҦGU,�oomU0C�C�|KX#o���n� =5�k����
(��B�6����Q x&���=�]���a����6����V�l�(e�Mmy� #z�M�3��U�kb�d�=��2��{�E쩶
��1�װ���.�����?0���9k����Ej��
>�S��2v8��b�7P�7͵b���$JZ����j�!�AJ.}�ɥª�N��OE@P�'`��&�Ne�@�b�g�L�T�uŊHT�0���#�1#���1C�����v�{k�~z��uơ���O6�cɑ�c߳-�5��=��)�c�9v�RN��,1b��XY����Z��G���Dl!����wdJ�o�����Zq�a�����bAiۧ{{ӕخ+/��I����R���X����}��)1��SK擆�ʏ�_L��� ��<QjH0�Y�U�� x��&XR��U	�G=��%��H��O����E����i�𻯥0�����B!��z�4*�i	o���j>��9.�@ˁy���T7��֕��������L|�X����8��1~J=Kc��/�e�~�5�;�#����$�U�}w'��^�#7<��&�"bK��\��k+����\i��x�0��n%��v���ǣ=8�F&;ۄ(]JEݶ���n�������?=%ɂ\����Y� }�d�+�qS��o�y���x�F��I z�c�y�=��3~Eքlc��f�ÍC�+i:j��6w1۶$#Ӓ�[+�/�+}��&or����rkx��H����y��ͣW�����t�"�6%�ᖤ$HYRt��̾�U/<�.e�8D �oSQ3�DWq���-�riZH�׵�㤚ʞ�!�#�0���K�R�uٮ�N�M���X�h����s�U��$�Z��pB��z��:�ǒX';��!������t�������x�*�u���a�/@���"��[�d%����1ҷ���:ֲ�J���z�l&�}#7��y��H5�tu��@��ֽ�u��E���O���X+D�K���������˴�:�r]��D�)�T���e]P]�pG�9�+5ё��Tw��^���<�$�r�U��	=u�+��Y�s��'���C��N����)J<�ˆ�氜D�/^��~��Q��Q�{1qIYGw|��N�z_ꃳ�{�w�<$O�"(Gw�Z>�x6"�p�I�������/����޳A��c-@��S< �@�E�^��l)��<��*e�f�L�0n[���kz����I�\ ȍ�?��]�(%�H#F�孱�ٖF�L#�I6�R�����nO�U�Z&;���;"9��ri�k�d��r�l8����S,&���K��ڔ����aɄ.�sRk(�Ffڔ����{�u7ހ��t��d�N��%%�t������ˁ6����ӵt+�-����U_�vq��5af�,�����]aE�_
?;�?���B���7M�;���ф ��K��Qs���'�oT�J��*���6\��/^9��bY��XV0|�p �:s�23Bò"�S�L�?S�ހ�߈&/~γۋ�	~9l� M�N�������` �$��b��d�N��Ud,U3�p��fC$X��o@����� �T��;��v8�'�v�^9������H��)���'���'�ß���]�����܌8�)?RD�R,�����TRZ��'7�ϥsi'&�����I��Tf�A���Y���x%]��y9E+���d�j��s@�-�9I5 �2��.CYԎz��!1PW��d�d�_\�D&E/����^w�w��M8Ә�d�d�W�gzȓ��.����q��{W�C�F7IW����5D����fs�I������
*o���ϥ�V���]r�L���Ĉ䃲�[�DĔ��ԷJYwf(��[hkK�;�,�=��GT웝�x�M�+|�]���T~fہ�.������{�}j�*(��!�{�L���:��lM/�4���U�&ol\��t=�>��zw���6�XLП���m,�<�L����i���I�i]��X��ޫEkd��!Jrl5�U�_�m�g�"o����exT�����^�ʫ����HN| ?��r&��0��h2c��_y�&���=`��7j�\k:0�� �FǴ�5�p}}}`�Z�������E��RL� 2Z`��u�tA��9�}�Ɯ�7���y(A�����)��k`�`/�|��� �v�k_qP�Ip�j�rO�o�I\��ٕ����i�*\�_!�A�����s�)�ec�W�'�wE�˱Jj�4`���8J�����*O���+F���=M���	�M{�
s�L��6Wu��hM�\��=�,�ƣ���OV@U�b]�n:[��S'��q�Vݽ88e�W���;��%]|i�w�9������Q>�����_�觑6��x�	��|����A���Y.ئ�2?e�x��T)���Z�8nlgU�3x��<�x1�(�=�@5�(8���/�[-=���d��K�s��O�����^���O�+�amQE�vUhr����6�\쪬%5L����;�m73�H�rd+_ ��H�� �B幦C�DZ#��tS���8���V��<v��iv��2�=��$���ଝϬ�>J���vTz~m�x�F�@~����D�2L;�Z�mo�x�a]�Ql��*	�?�b�"5�F~���-�����,�p "4���$Q:��"��|k��xfW��/n3���=�l=�i>��}S"C�2��G��B�a �����=��C�2yd�����x�{��� P�?�Y�>uM�ע�?M��4���T�HհKFf|�R���!��ߋ]�w�%'��`�P~�cdw���;"�����G�}H�U��C;�6�����P 6����@�	�9��o�PCIC�m*�rP|�t��7'�S� h�
������א�����D4fO�%V��OJz��o��Hh�	-�������C��yl_F�~�^�S���Hz��k�_B9�O}������l��9�/Y'_t�R�:޷5�͢���!����;y�^����59O����n��n��\u��˽۸�2$#'�>W`LBw���;L��.Qg�j��A�f�1]����~�"�cA�w����W�R�k�՚��j�H�����l.	�:�s��~=���@��dI�i	-�4�A��G|ӜP��'()�C�Bf}듎�?�h���ڟ�?�'>�yW����,�8b�p���]�/�kT�I0r�����ɬ~�F��{��DO*���M���]�M�ݳ)��g�czC��J��r��H6����,t����Īw�O�Dm/����,�KN�47o؟���T5&n�u^���VW� p-���S�p9�|j3mp�Tɳ���v�,L\����q�"}N��V��N%ۀ��C���қ$����-"	���7l�����Th�h�Ⱦ��r��$�1H�$̶N�aB�xz�ߊ��د��3�B0�h:�39��dS��$:��T&�����*F�V�j�le�|Lt���J��7���|	ҞUMLɱ���ڶ�+�9��x���3��\ܳvL����a{���n��������Rl�u��'��mʂo߳�̛y��2V�T��$��y�T��<6�LSz�h�hɃL3_pP��N��kW�M�g��v��Ȑ ���l�3��7��L�Lao��p��ޙ��ǧ�B�V?��Yw_n&$O��p5wО�K~�n�-�����{��_������2΍=b����6��=�)"{J	��K���5T&v����֪�^4ן>ƣ����=C���q��z�w�@6l�'�DG�doR��s'fߘ�W�I��=gK��:
h�J�k(��Q������W���<C�z�<_�m�����+�B�Ӂwȅ�{*췋24#If���4 �N���*�t��85�5:���N��6�PMDR�7����P���*�N�X�aC��WMM��ݍ�Tv����'V)Qe����N�D[`ŞF��`�aJ`���i	O���M��u�cP��E�&��+b��K �����F��Y]�^B�[���L�����󌺽m̠���qN7�V�dq��2p�ڏ&�������a���9Ÿ+���;54Í���>�!|��0xo�@�}�2<�'i�O�=��/D��<'J�E�����,�~i��I�:|<}*�Ϝf�����XK0|2�TW��q3!e�����gZ�-�;�A�M7�`���9`#��"o���dݧz�ꁈ�����A�H%#��O�fw��_������t� >��[�R���M��,V�g~�o�6`VVVB��ru���Hˌ:�O��lU���|���Ae z÷"y2ٿ�<�%�H0:ڪ��iR�JBUpqө��j�y�\���������,�ϗA[:���F�H�{��*��)�ß�ͤ)?�5��E��C�;cd�0	��eG�Ym7� ����)N���'#?��{k
I�-N��;�`*꽧��ݢ�x�l5KI���/��w�oG����LΆ?&[�x`]g������R:����Sǀ"㳣*-�)�Q���;O0�����zf���{J��U�vr>�G,6[���]F#!p�d2%B���z�	�9	�2����'��ޓ�,u�}&�s�ې����dfe�<�5'&N���9SJlp�P����NE�%�[9(����m�a�w+X�x�<�g��g�<�x���b0�\�t�����P�tg0;^�a�,�p�OJ���|ܤ�{����l���,=9�t�b����Q0�1�m_���8X}=&�������	+��\�2�!�ɉhbX|�n�}M�=e� �,�T����a����mg����ƫ�P�@ 9�J�'?!G��f5Q�탱�?{��_<jN	�O�Hm=V�R���*��[��o��VU {j�2��O��H��x(����k��'���ַp:������K{1>�~(����u�b$M�b2.V���q�' �t��v	W��ƾ,�;[G�%k����D�E�H��rK#o����^rN����~Pq��i*���FQo����,ۄ&XL����+�`SlK�@s��|p�{�{�ʇ�B��;&��_��>��ۂ�hߔMK������W���@��Ģdq�#���<�/߬�:�G���Q�����%NvF֢x1�$j�������S\zڵ��	Qz�?3��\�r�}+D��6�r���T(�?v�)I}��+{�W���+�����?���D=�,�!xYQ��2�[ނ�NK��E+\md�c�[��n=$QP�Bsb��v���`Ep�����8n����l�N�o\���[�B�� $�f�}G� V�U�R���GH!x�&�l�(u�+{�2W�����)�]@#8����~dx?tJ�1��%F�
-y�[����Pz���`�s?�6�J�K�����Ƌ9%�`|�">'��j��ő�>X��%�޽>23��$������q5y�qC�t�������O�^�ۓ�}��H�1i�Z��h�4��м�K?�b�F��E�9�+��Te���g�N0���ܹ�U勉BcC��B$Y�B��۟/���|�6�2v^+i��
��r|C�X�Sά� ùqA�H<?{xT�^P� C�c;�L��P�V<��EMN��J�w���bf��[d9Z�����]6��n�#aΏ�����R�J �Z������n��ӫ�@����MN��p��L�8?�I��������ɤh*�`�g���[Z��U�n��?���j"��4^�Aq߹�<���}�"NH�zF�\����	2m�<��ه4��h%?�`YI�=��(�Z���9�����>�<ݿ��@v�����$���DE�ư�&Ss�`z[�1����x�a��0��`5>־_�헆%�`e/�2�]b��߳��R/��V�&*��d<���/4��}���'t9ҥ������}��o5�o�3䭒�� t@��y��5�;>%�g�"��c� k�s2Y�=Jv�{�Vq�dP����<�'��3v;�Ǩ��09,+a�m��,  G���iN)��yﳛ$*�!�̠@@�Q]Ϧ3#�U���*�$b��A�*'���өs�k��k��uU�k���97v�9@��B2粰���٢�K8r����[Ò�h��!@�WK^��������g?Ϧx�V"�e|t'�ڵ_}�%۔����y���J7������VW�*RJ��x�7#r]�q⪪TsO�qU`�������/����f������ITM|w8<X0B#K!� �şup
 �����XY��ԧ��X0�ԙ,("�>�$���s@�95�&�_e�Џ�9���;�w��r�[�K�B�Aۏ��������k������owC�����@$ň��L%u�Q�r+ƊSU���Η�D�� X׵ՒC�?T4�
���KVy�ާ�94�x_����h~Y�m�h��&`�gR����yY-"Z�YN�����\��K�)Ù4���xL���s.%7$!��G D� Uy���81�����0^���<�u�^uA��/���oPa'���ER�9W��ts](�Ǔ�C�]:��li�?5g��m�8����LEUD H��w&�D䰋ML3wm4�s~6�����ƃ7����m�<��Hi^�"�@��hVT�9�&�|�>�-Ykٔ�#�dNPn�iN)BaD���1b>n�]&�w����}�nV���=�t�*��H�
glTͽ��7��e0W ����Q�ѩ���z���d2��[U�;5����l�ˍo:a���,��Alp���,�1�-P��3��N)vݦi��i��Jq	*�C�'��S۷yG��5��anwx�f��"�B��r�׷�y�
��n>?UU���u8���l��BE�|�Z!"3"�p�j�*;yyr~~��X�"DT�:�WA�n �� T ɲ����b���c���U0K�y=\�-��xC-*3D�TM/���@� ��� ���{"���m�q���J����.��b'���!q��!� ��"u�j�v�Uu��9�~k�o�z3j�0K��F>�l,t���a�������dNs�B�	I�_o@t ��`�]�v�X
?3���_n����BȘY�*�ȅC\4�2|0D ��1*
K�4Γsn�l ���`<]\\&N��<L�7-݇K݀���J1��ic�3��e�s�B���d2Цm��"Vu�]X/�"R׵� �P@׶�B���f�U5�G]י_�*dN�Z�5"����1���mU�yod�{�������w�lL�kgd�<w}�*�p�~������%"���v�Λ�<0Pf,L��OT���ca+�SնmS�Z��+�� y�ez�����e�`@�H���A5�D��A����1FD@��>"xG&��%��iZ���������\.��jE����ż]Y,<��������A;L�o����k�?������q�n�xG���%,y1�LRr�N�L� �s�`���Հ��hT�5Z5R!�����ttα�|�����������۫�zT�m�um7������������g�SA��[)p&$�]���ߐ(�3\6c9U@cE�+�$� 3c���ªe��7a\/6o�?P�!���J�T��;��E���[GĜa��Qx�� Y .B�k����ۑ�, "�lA��Z-N�� �̮���EUsU{?�繗l&�Lп��d�2#yD��A��� ��="9W�����<� ������Q����k��w��hk��?�06��G^nekJt� �5�*(7l�������=�a��B�j���D��<"Ɣ$%Q0����)��M�}ЖBg��;�����0:������Y�|������ߥ��2P	��ǣz<�L�ە�T!X��"�΋���n߾u�D���PE�'GJ�9|�Rc�Z�'�mK0՟�f�(�Q�CVۆ�P��c���6VSU�2��:��*Q��z�DoZ�fX �a	��V����|�P��ϒ_b)��\A��5ZD,�QH@D��l<�X[a�u�Hs�2�>v�3��z�>9=}��w���.�/�����G 2������|� ��C��޽
�g]�ݾ};���_���������/����޽{����˓�����s��b�x���l6��~���_휿�V�ɓ�M�ܹ{����W����QU�}ke�7�7�����m�3��wt͑@sXm���O��x�����k�ۮcΠ��uf`��|��RR��x<��تzEX��e����c_���@&�g�a~n��/�:r��CGP*� MZ�HL�����` Z�k��P�]Z��_C��H�V�j:����a��;en;#��W����SJüG�{,}�U�o7�]��I�"�������&���@�RK�[�#����X�_Ed�Z{r5��	T��Оl�B۶���:�#@�.�$��> ��������V�����aJ�m rU��z�޼<y�E�pˤgfQ�������͸�s[�sK�`�!΁�
�,{g�s���:�!@��u������ײ�$y��2'?��&�q�	[�d�ՌA�Ӌ�,��͍¬�,o�~���!��g$t�����!�bF�}�W����N3sbU�1�Y7;�'�`ą���W"˕Կz����.F�t��Y]p)�Ѹs�}<gA�AG���WA�K��� �Q�Y([YUMTr���S���,�a��(]�%x岍g)���yH1ڻLk��.���{I-#�����k�HU[7R��J�v{ç�����vaND��p*�~�oAD�<6��r����\�W)t��d��v�Oga3w�� ��2���\�׋��|zM����DeQ�R�w�4�m5#����m����
 �{�Q�a8V�)���o,o�� 
`�ox�� �^��&������p�&�1s4Ŭ�����+d���@*I!��f��b�Y����2��

���0WU��P�|��֭[��t:��-�^� B�]ׅ������!���Ȓ\�Q�)v��m��m�+��:�d�9!h��{o��u]h�˾�G�`�̡�ƣ���%W�j��:��� X�1YuK^	}�V����'�7n^�e�6�{{{U��Tă���K����TSJ�YR��K���s ��]�:כּ���}�f���ݼ��2�����R�ӡͼ��gxU�<j;���&)�9��X`.,����)� �sѕRs�B(�a�H�%"���
� �\��G�H�-{d:��WT1�Zr����bFz�P���J���m5Dp7�]�����Tx����p+!�,�m��B5�G!���N, 
JU�ƣ��%��3)b�r�2'�Ս���{�Ř�.�`"1ƮkC�vD���1@�EJ�r)�u�:;eJ��M�A�y�E�Y��<n���	{z��Gs�n+��{�g�]@���	�����**M�������
r�N��i�*t�T�|��}�E|���*lP���BD  f²��u�����D.�sֺ��]���z-"uU�����&ha2����|�sx>�;_�o�,W�h�>��h<�����`�S>e�x=j��ʉ� �j>��$	�Qv��B�����>��
P���˦ ���^���B�~�]U]�q.]A р[��4H=En�̺=��5�6�D+��{�g-�`�nv��ΰKPX�cfP G��{/Eo<��|���]a���@߬�0��7�&�طe�v�,� �����Abn�f<�����m�u�(�D���^`kJ��v���J�k��`iC�ko���y����Uި��: =j�ðD�,�x��XehF(@z7�֕s4�R��jm��/���i��6�D�\.���<x0�MMG���1�2�y�UU��ŅU�pN���c��Y�qeU&YS45a�bl���cLM�i�61WD��4��i��ؾθ�}*m�ܼ>K7Z�r�'�[+��T���dS_�B̬�q�J݄�|�]��̼ �ΏF��dBhg�!�snKM�i;���)�Yk"*�m"�RL}]v��Ȏ�.��-X�v����4��}��p��Ps��wbVG��tQ��E��  /�^��G5���nfEt��.u��l�N�#���9��,V
�	r��*�3o����~����N��s�� T,�A �|��G�BE��>m�Y��k,�<�T�J������քU>9��LۍQ5Ip.ƮmSUՈ�G%4'� !`�SB9�^�v��ք艪�&r,� EՒ�P�r�s� �<y�TY��"x����u�����8�٤�"�)%_ƪ�W����1�n4j���2ey�XU&�*h��5��ȁ"gU"P��3گ�ޯ�P�>v��� ���_on��̨��6���4��΍a���+"���ͦ�b�ҶQ���8g
�(\4��"d���nb�4��EYDY� �3�C�]�)��[oEU���Q����5�<���%_=�wW]�H���i��՝YԨYt���h%^�bfLO~��W���S��������d�m-($��k�&�n:o�zجx?�,�y9Ղ�eD�0m�]��}����$ ���X�o��f�Dz���������sΓG��r����gϞًb�2��fS�|ہ�:��ۇ������N�x6QZ0~���)��%0ھ�s��-��z=N������R/����R D�s.q�ڽ�1ủT���M"K��K�4�m �Ȫ4Iх@HM��JW����������*6���")%a�ꫯV�UbvΩ�Ng���|��_>�Ho���d29�8�o�q��ˋ����|�{���� �޽������_<}������w�===}�������o��4�'OF��ÇG����*��p���7��<��v`ggel0˹#�.��7�2�5pHР�b=�C��u�j�����z�i^D�B諺Юi�ؚf�����ضV�L�Axh͜�o�������ۢ��7^�ʌK����~۫߬�)���+_!׬�z&'V��Ek �}7׺eڹiIQ�kDD +����^N�l~��2Гm%@�G�.�06/N���y?t�b���j$��H�[�
��� ,C���#T����NgU��ڪ��ĝ���ȍF#�4k��@Y��Y�zYt=�Q-�k��Hh݉M<��k��x�΋��J6@V�%b�D���K�(�TQ$���s��.Ӛ�˨j��`�]��br3�-��z�9û�'����g��o�jUT����^��H���x�]p��+ne�˸6@���%G��9S�
!X�8̪@7��6�Y~����bR�'��������	}�Um�b�s�G�L"�ݨ1%eaNJ4���Y�4]�zD��!Y4�7L���l�ɔ�s�V�vC�����ev���?����m�����^�0��{[o"V�����C,� ȹ�W��.�?�8��jVt���G ��q����q�U�}~J�f��K�9����C49�k�,�r"
��뺮뚊^:�
'm �ؕJΏǓ{��`�qoo�9wyy�R��*[�e�f�p���s�!7�����Q��lc^��K���>���-I�����d�ҵm��ͺ�z��	n�(U���xT�5sjڶ�:D�୭A ���\�v�\ݺ5�MW�Uj�5�r��ID��
UW�[���h��{�S���ψ�燷o��կ~�l�����}��;��|����������'O�<~�������4�'�|�;��;��?�?����>��֭[������������/�菼�=�b;��(R�H���d��1�� b�bYpLY�B
�_T�~[�
v�3DDrb�ʮa������Z���4	����f��mБ�L&��؈�)&��L�p��\�����7>�o1�����?`p��S"S�R;�o�ޢ&k����[�*��Y�C� J
	� d*�I���lͥ�Խ{f���-�ד8xZ|5*��$@�yӥ%�����Ę�D̅PMc���VדL�EA�M/<vݦm7U�CJ���j�T��TUMm�:�T5Jda R����D��ʹ�������E�QQpd{Z�Y,�]Ԝ��]'̎���"��vL��0�s���$�D��:k�cK�Q���v�-���������v���%Ý���%�ma�@b���"��.�>�����cJ(@�;@���#�.�g�2�r�͙�P��)�����[1y&Fel�|�m�'[j	��m���HJQDY�t`n��9X/_n�Pcl�RR�#�(��l��ɯ�>�sS�`f-��6�n�RT>A����n5K�H*���G�e�d-|̜�� �~`���hjĲ��,4���o�7��cK\X)+v�MiY������n�댶�T\�||h��m������0�e��q)�2�����,��ش�y'�x��0�݉�Z�����鉉S���i��v��B25;�;�J?��48ÇzՇ�q5�Uj:�6�"�H�@D���Ppt�+����t���[��w_^�I��[Ȏ؇R "��,T{{{"���4��L�W5*$ �����9��]]^ߺupxxu5o�f�uU]�bB� �ؽ��[��?��/������j�f��jյ�TUB�b��cN]��������97�B������'��t:eN������I�4mV̡8dj&:��\^dġ@��� L�
Cf�AV-^Jɺ<K�	�i��&=�X� RJ��*���1f���USaN)�����bJm�2�j�e9g� C�a��؟J��Wo�zx^�k㈈ h%��3uF $��Y�㰩zB��Lr�䟋�J��)��[���l=�]߁�6N1�b�9[�;��������^v������5ܤ�W̲6"]�l#�	u�h��u�;S��V �-��V��D�Q��po�[���$�n(�7ʻ�%�)�H┽IUk���q+ݏ ۍ� ��ʢ"���<��f]�Ց�옡��Z��0ǘ:N�vkiť�����pB�s���G�D�u4����u)�d�+D�P����2T:��oS��=��'F@��ݸ93��a���6��՚����8�	��̕!�Y���N��h�C��`��Z��J,��d<�Q]��0sJ�^���*8�wɊLɪ��&��I 	��E,�d��n�|����KY��&
�~�5���΃���8��hM�m�s���|�%I�*�P���2��z3���T��n�һ�Ka��j[E=�� ��˱�*�λrP*�*j�i_��^r�FX�!1)o�u��<�I�V�j���,v�h4Z�V�oEa�]�PM PQ��jd~o��O�ͥ�� �e�:@1��_%ھ�O �eU|�܂Lr�or(�Ȧ�`�\�Mo�^�MM��u��O���
m�Y�$D��;a.6�2  5+duo��V����d63�ZU�e�q-=��y��{�}��"�ٟ�?}����zr̼�l~��BX��)����O?������G}tv~~uy��?Z-W/^�`�_��,�Y.��W���?�q�i۶m������.����w�����d�k;���Ήn�w�l�Q(��g�� �BQ(�G.�p�5��Bvf�"u-16�JJ(*��h4���[G+B���>KQ� hc��y�4>�����q�Lt�H��u�B[��	6���
��MW�%���pf-�|�]�O�m�ٮ�}��G�V�q��Z�Oq�r�s��}��크j�Bp{0!d('�_��W���5��:��+'L3h�S�U�c�yD��U!pJ]w�;�Np��*��B~f�� ���E8�Fs�m��C9$>���>�煄��Ř�uU�UMH,l��4�\u��M��Y ��� "}�H��m*� VƈJ�!� ���"�E�M=�ż|5N��9&���cU57�E� ��"B�MJ��D3A����|�JV]�����A�ˢw'�������L�0y��,�>��@�1��,�C�ڿޢ���M�!�fy�, ���-�麶ib���mץ��>�"�Q\__�۽=�	P$�k1OoD�y:|�>{��oq�y�*�@@����헵� ���IF:
ڶ?��� Ü��Q�8�0ps�)%N�o���<��i+�
����m;��sM�7o��$aU�U �@�։��n\L���"�j�z��C�6m�lD!Ʈ�C�qğ�!�'�s��$�\�����<A���u�`����P�R߰�v�����A�`i�o:1�;���lٛ7�k>��Yeuˁ�4y���l朋]�RR@�=�
�'��*�>� �����/�����tv5�+@L� �S�g��Ç�o�.�/>����>���_1��b����/�#D��>��;�sΝ_\�G��ŗO�>жm�={vzzf?yB��p��g�;*�b��2#��ܖ8e%S�S4�4({�	5�V���a�΂�L
����E �|j_V��6aj�4�b������um� ����ڶ�3�9�X7�i�ylx���SrD&-�I���(c+��Mё��p�k0t�Į�܉B�R|ӕ�b��e:���+:��6yP4�_b�f�n:�UU@IA8��ATG7������DZ���a>цw��O�s���H����
���ڳat�	3�VU5��wڵ����B "K�i�od
1׬�s��rkFIKO;���KD2b�[�V�o�c�10f=r꓊�����V�l����Z4��L¢�n��=_*;�D��5'$O�)��;�ܖ}#jQ�P�#W�ľ��#�f�f��#r� ���2MՄ��t�p� @(����r#e���ͩI*V�^һ ���$��3/"�ΦUU~h�Hѵݪ�Δ8sO�lC��oED��w���{H�F�W��9�D���u�B�E!̦���,���;�u|L�5�FUC��J8���'��!�Ff��4���t��i�����o�Y�o�G5 �  z���Mܻ�G�?��]+�������U��7_=1��ϳ]�g�E��h36��UK%�"Uu�C�!�'cu�9R����Ѫ��\UUu=><<9����������R�s���}�Q���CE�Y�|�H}7 ���RUN���r��Fj�ɩ�(V@�}�:J�>t�M��8@�d%�=0�(�k��lz���"�?�b{���:x��7��i���@����W����ݥ4_��tw��/.~�������z�:�8_��1��|���P��
�����n9Z�J���K)dZ�i5X�`G�9�Zjw���h�5���N��W	O�N��"��V��"F��W���p�u��d��ۢ��i8M/*>�o߾}����juvvv�Ν�l�����r	 >x����,Gt�գz2�Tuu��ݦi��Yg�2r@؇)v
n���̉�������D���nx�A���R���n��4�����M&s! �������2U�b�G �r�f ɝ�o�Dj�Qf˴�f���٥����N
����1(����/��H� B���V��.�A�%��L�����^��i��o]?e�ؙ�J�m�̵�rJ}���i�嬴ָV�iM�X�v(�a�l�s�a	���$Ke�gΙ�����֗j`aK��~�
�c�y"�p�`�S�Cp6����U�M�r� @.���y�E���%�R�$�T�B0
Qs�Ma��@�?��.xfN1�F#�b��#J����@�Xq�eJ>n=0"��EeP���(��B�ƶ(���`���~:ۻ����ڮmb�\,��*�,���^C��-'�D�a�3�>��1�^;ݯ���[>y�5���s�2��HU1�P�_��Yi @$B�i����,W�����7��w�^7z�+�q2q%ڦ¯�+���&\��/^��]c��9�b�! :R͚�� �������\D�n��o6�i3��ʳ橔�?���c9���Lz*��$�h�"��#���r����D
f��""��'��P8������1M�Vw�j��-�OV��ps��#�����noo/T�b�X�7�*d��Gn?��ǜ�VG��f����<::���[.& �K�9�_���W��s��l���'64ˑf�UM��yb{~�s�پ�9�:�B%B�=��2  �>���2� �h��� � �+2��kp4��B9t����̣���������J�1*�I���������SL��\DR�mۦ�ڮ�r��u���N����U�CUU*�l�"X�k�uD$��/��۔�o��;HO^cp�Ôgf�2eDRC��Ҵ�[�����&i2��Zm�����_�ɓwR8��{6�Z%[��-���o� ="8�`��JO,K��˫��7�(�	�Ge_9���hx�/%��W�B�*T"2��f�Y]�D���C����"榛�^۶��U]��c���'�;��V�ҼR����!Oby2� -r.����>/��W�	f�� �iw?fd��"�:f5�$�� ��U��&NWɵ�[�����S-X  ��wy=�aqދh�"yae(�b����ì��Ptdh�0��sTa��R��]�Rڒ=��a#���m%[���G��Sb>=;�G�?x�����H(�1F�]]�֏	�9P�&�5
��`�e>�l�+�-(��m�����O?���E���_���#猔�
@�/������f��j>w�&Ӊ �Bl:p�'�1����$���Jm����7���=�,��o�'�l17ph�ˮ�\-Zͪ�*��&e��& ��υ�5�ټ�	{��lx!�f��l����vG���N&�zTo6�����!rU�G���!�4�L���e��k�.�X�0��f����~�)��C���;�'�=i�k��X��j����""�'�L8ܡ��	��I�F#;΍P�V�V:�C��Ƶ���jVУzDD���Z�{k�������;�O%1���u��k��F�U3�.�j����R۶������Rn	�����T�}En�6g�g��G�����۶i�������|~vzj-"���1���$*,�#��2"���Ƙ���Y
$�L��Y��|f�f��O�D��Q�-Pr9#�Ex.���J�h��!	���Q�OScC���	;��v6�%*�\]�W�ˋ�U|��>��k)��"DO��G.��Z���g�8]ͯ&�I۶'''�%d2��0qa=) ����ys�������,[��\"�6*��n�ٵ@	�e�Յ%ӺE�l�-�ը?v�.Dp��Л`��"L�L��A��\� iE@@T%�Ք�%yEHPn]�!�^.榋ȺIh۵����
��r��Ap2�<�,qR $D1�0'�!����9��lQ�11��k"��oۜ@�8<p��됶��� �k夠`u�,S��:�j�lRL�Ȏ���nS�R�!zs(�c��l�rFѦ(�m�{؊��;!���|��_E���#V�OIbdӿ�W��-8�}yg�",B�y
 br8�\i�0LLgsL���)�n�=�z�d�m��������><:<���0:���b�i����9�b��Ɣ�[z��@ ,z89z������}��*TUUוv�9G�Ω�wNE���j�3��]���3�4O:ꋅ�T���kR�k��}�~^��?M�:{Ԥ����
�6���*�nݎ�|����]j�vN�cV�׫��N���d����l9s�*�=N J�v�?� V�~e���c�@T��af�p�>����|U����xu9_.u]M�Ӻ����W�ˮ���(�~��_%���w��2�:F}5ڼ8p�wU%G� *C��>�X�&��2����U�}T���,��li@��)� 
���"9��ܢ)7���b�$|#�c�~_A��=G��7���Z�,c����M&�\J-s�(Yy�h�䤼ųfǚJ0X/���燇�{ _ C3q��c�H�r;�z�yAUaUP��TY�G��ꈤ�s�15蟷��vֶEk�����}��fq�WG�X�]6[�������/�f_ ���K�n��I8W�"!'^��t2�N����68��&�����x��/_�|����8��N�D���ҫ��Dz�$-@'l�����1�Ū�hjq�����!W�H�u��L?0�[����#���m.͙�|��l�}�w{���!�pL�4>����g*#O�-��[�o�-US�Юk?��# M���O?�n<��ә��%*sUW�JB��>��ٳg�x���d��R�B���B�2��!+ܩ1d�^�#��̢��(���B=��E;ϟ=_.�U�'���f������7w�G�����*�)ߤ���S> ,cȨ�Ͽ~��������кAY�u�HPH�@K�S�e�y�5{�(��Z:�f�U����۽s��XKO��Z���30�WW	""`J����Hx||���g�����//�'''����k$$&UΑ& }[���ƌ�^s�����#ɼ��K�$?�,uλÃ��RJ���;���q��뗃q؍M����j{�p�1�m��~�zlr{xoK���n�׍���R���ﴱ��(�����L�~p�����ܻ��wt+_q����	����pE^)����
`cBDu�%��&4�ƚ����ڪD�1stƹ��9u1����әa���HƩO)�Ywg�{y ��<�z�S�d�t�T��џR�ëw�ͣ%G�\�6m��ݻ�y����$�^r�9�"��@��(�3�띷DRJQU����j�PP��f�O$Fr6�a��]��G�Wד�x4�Ȧi�a�v�m�@�h����������痗{���ѡm�.F�D�x�]ס���bh�L��w�A�9s�X��&'�;���b"��2*.x�nc��w��b������,~Fr��kø�7�Kߋ2��7�HF�PU��]59���{�u�z�� ̖�k�V��F�Ѹ�Z)�U/a�$m��o�Wݝ��+�E���%ր�~�����x���.yF+��@�^�����U��m���)%罅��E�m�k��o�o����Z4��Q�$�B3��"rt0���}`>Tu�Z��P۴m�U�Up�3G �UU�s���K�\-��g��j=9GjD�7l�0��w�X�n��U��{$"`����$�B�f{{o��F]U"R�������//��5�����
���S����_��'%V��`�v�7��"U5��ɿRfJ=<��(�����s��
�:Q@D��)��BV�,H JYX� ��;ƚE��g����JV[�ro�\Zc! c���e� �y�03���ɓ��S＂N��;w��n����m��k��R��6�����ǆ9���_e�F,�h�ص-�FjY�
��o��������m�h�xxHD^ͽ��n��0���B�C��{NZ�x�%��c��J�m��[�z񙵀��A��������C�FWQDA%�����L+�1Khz��8�ƺ�a�#",؊%�˱��'Za��mB����WO���OC@�*�8p��9���-@TA�@VR����<�!殦WWW��"D�(=D@�w>q�����]C���6�oF���l�]v�%"z�I,]"��,fG<�w������&����*vq�و�����߾u�b�:S��z<���狗'/W˕A��ITW�姟~���c�٬�OK�O��,�v�!���H�E��s޳H��tm{-����6�5��m�asꜰ���m�����e���ݼ���CG$�R�i]О�dW�U�R��P�����'�Y�s~�Ȕ: 4�3ό�"����@�����چ��`l�w�`mU�hC�ʘJ�������QW3�T��ZUmۖ��+	 MӜ�����$����y/�6�Y��^-���Z�^kǑ�p���i)�����8�9����G� (	1�F{�r�P�0r��",�51W� �ʁ�l����C�r��D�r+o�����)����;�qq�_=�M 1��F"��*B�Qq���_{��� �#�'n:��u�
w�(�PV�Γs��* ��.�d2�������yv�"�A6��Rn}������ˇ��_�u�7����Msrrc��z�X.���ۖ6vf��͢Ȁ��;(�!�H���e��z��c��� HY���VҖ9/0*1�B�u��ūUة�DU ,���v7e�Ɂ*	�&��;<ƙ�R��"���s�1���!X�W��`n�7����$���m;�l���.8��w�V�'O��ܟȑ���[MW,��*P��f�ncJ���G0�;����妴�lQ�u����;;Aw�����䶻���+i���ˇ���M��D�l��H�X���r�\t܇�b�9��p�k�U��/�[�P�ɨHD��H(h�B�jX١�mƼ�P�Ӫ.�9P$7Y��_s2�IН&"�/$��w�
���"r�2ed�9�!�2 ƔT�P2�1%D�P�U���<	U�[q�p��U�!�%
v�5�-�B���zt������O������N&m۶�f<���ƃ۷n��'O�e���t:��Ճ�r������G�5��9��fGG��󮈼|�2��WR%��ЫS���z�7ƄY�SKn���ԡO��&DN�E�٪�n�z��ع�#aJi�X����u�Z����u��u.W�Q�Χ���.���� Yy����	�%�����,�`o�*��~%����E�|]lV<OC} 	���_	t���uM�UD�7�V��� ����"���,1g9��8W�$Ѩ���}�	���7�y����T�Vf�\���U����y���	7��
@Ű�^:��\5s&ܐC���qN�݌٢��Hbq���V��(��j�s��^�iÒ,,��m�d�.D-Q.l�d�������>�6���"����ċ����f���\U�}5�:$�|�do�8�=HA��@!�S�rCi[���II��2bxtt��o�����z�X��� �suRFBx����4�r� ʂͪ*ʂ����׀&��������J[�TJ�&v��Zղ�E)\�1pD�2����e��*�\1F��_�6�
*��@�K<Y���[@�:���֚O�y�V\+}�#��ɿ�"�kF�������M��㏝w��ݛ���ż
���~�Kq��g�wfSU5�%F�3م���B; ab����@����ך-p���UȌT��ܰ
Ln�~O�]ٍَ�s�-m���� 9 ea�"%)KN�TE8�&#�lY�jX��'�=�\:Ov,	��lg� �z06v�9o�A�}P�"뺪�w��T�nF��9�=N��������܎�؜�R�Y��薩��2��b�Z_T�����l�^��wQN�m5 g���5$v���t{{oq��O��$q0�6����������f��ǿ�{����~�ӧO��ͦ��[��>}�t���>>8<�'�����''�u]߽{����{����9�8'193�p8^�k.i�M���? d?� $��N�y#� ��mmשj�>�%e�-~���ٿ�ܧ��e�g�\�V��x✋1"�Qr�3@�������r�5 �D53����/ n��v� s��S�������]HbY3o�a;G���a�zTD���.�Q4t�˛��bd �N):�U�ȥ�D���(l�B�z���a5g��b�G��mTѻ Y���2�B�����^�7�	�R��1��O� �
y�"F� �p7���Ѭ�
�*F�t@*m��"[�Q�b�]l��eTA)�\�.�t ����],ϵ�d�4�ex5���~����� !������!a�bK)�j���" �B]tYJ<JDD�R2�
��P�a{.t\<��6���Ǔ�[o���4}��b1��,} f��ёGX�����#�Z�u�C�b>��2j��,xi�z&q�fU���R? ��y�ɠ+���K�E�)xO�IP,`�AkR���͌�L�jX_��� �2� �C+3�����5FО@�򓶅i6�6����o���ݻw.�.s��w����ב 3�e1SoIUs]Ʌ�����m���~23KJ�tG�ЀH�7�+�m�͠i𪕆�o��缃�h2f�v��9K#�����kj�v�4�
q,�uT����GI�t��@Z�c �RRI�N�IwJ|@:�SPb4Hi����9z���w~�gl��{���|<��}�R�s�"����/(�s����S���㳻""�(�� �A$�����j��O���N(Pu0U������"� 2 '��W8U�� ��'����7I$V��ͣ)l_��&+�2� ���#H��wR�8���\��Iϴ�w�0��<
g�	C�r>~�P�W��f.��e���N��t�p�QG���K:��V鮶����RIyl{�:a���唭��,/W��7']�1��=����)yI�F�>j }J肹6(}tˣ�nLi���?>��L@����/�)�I*(���m����4��ϥ�O��.�Hh�TME��6�3y�"Q�_�����7���8OO�_�"-C�� ����,Ѣ�B2��+�_vZ�>uc24Q���t��iL!yj`�{��JΔ�������� �_�������h@��"��8���e�aQ#���q��*9}���������b<�sW
~�1�>L��<ܤ["�r�y�{�La��|��t*��L_/�=�u�VϝW�pr!~�pެ��4W _�Ct��(��5�N?1�x�������
�����8��{�����������fsu�U���ޏm	�7)�&���g	h�[|�y��'����厧S��xH�-�J1RyJ[�Ũ���=�O���hh�;����12t �կr{u��m������98���5�sɱJ~��jzL*#q��C `��K��"���X��C���\��j4���|䧋�.q���}2�Lh�8�(s� ���NtA�����n4�`	?���)��q���k�rɿ3���SR{�Ϫ+��2#���|m |�*�E@?|��\{3vMV�(�|���`�f5g�������Q��e'|�XPڀ�zrvp����N��F��Oj�>���z29�J���mm�]73NgE�璖�dD�!��O���x�V��I�n�w��#���e���0Ў����1F�hOѺ|. =d��]�[�,]j�K��lO���*h������q��s>�3�7�
_�ż�c��y	Y���%��=n���y��(����bj(�M
W��)Vf0���&ư�ӷ|H���ӱIohi7�����awXX�<_���J�<�W,8����B��v5E���,��c�'�g�R�i��x�f#g�u�<D�__v���[����?�.�Z��4�s���s�z�Š90�y'U����B��[jw�\5��*-�����}s��kw&F��k&(���f����XS��V3T}!Z��i��5�` S��`k���._R21u��8�SV���s�XVũ��_�I��U��Ҕ�cղ�(&u�~g�i:�轚�[>Νj�ɜ�o������aC�Fl>B,[Q]�Okt5 ��phz���A�f��k9���lTT���y��Gy����7V��(��Vq������ݪ�G�TP
r�ꁟ]�("lȒ����w�UC_m�){իF���"�`�b���/<�v
t���䌴T��r��)&~�������_X��	:�m����䙼�oL�QP/a^Sl��jq�2IT��YH�8`����pH�}F�n#gd�y��#�t]! ���>D;I/k >�� �����|��cì�}T��zڼ�����*Y�Pq����x3[�wۙH�6�Ε��I+Mh�j��~ҧʴ�E0-�}���d�Vcy����~�P@�p����_�D$.ZO��W�� ��%l�9�?����&>���XrgU�������Lۓު�"��X!����$���D�b
�z���)��;�;��(: c��0���-�6*ۿ,;�����.�#6}Lc�
����^�m��h�}���)a�Ħ�G��G�1�=��;��*���ӗ��P�(��}< �?�������6H'�"ֵ�d�7�Dd�G���=D��U}�vG_ϝ�AY�HR%�UX�k���

l����U���3��C�<��$�*O|��qٳڕ����/,(�@TܝX�
����;�>ho��8�8�(
�E�U�<Ԝe�6��|_^,�m>:��6?z�dI��z�z�)�����Î�w�u4%�(Ǉ.�
.ڧg��{?���	7>�3DUU�"C<l_�'��^���Q��I5�D?He�WGƁ?�|��K�Z�h�ݗqv���ӥ��x����O�/A��~���r��)��6~�T�\W
U�b�ʄ6&�������z���d+�o�y��F2Ȣw�V�%O�\];��AW������Jv��1#0���"����,��Bw�3>YɞJ�h�2q�[�_���~趠xA#t�i.��p AH�L��]Ndp��a�ji{$��˻����k�l�s���J�8�n
}�E�:����<'��5����zy��(��tus�bo^�C��nr-�H�X��pJ��3�H���>��zi�`���ɧD+P��B��C>[��Ax�N{-Qz�B�r����>�h'�`<(pE�gı�>@f�;�tIh�C)5�R��׳ w&��^Y.�ͷt[�Wf�����`�#��P�T>~ER��W�������W߁]J�:����Wa͜��!
i��˃�%��B�N�R��x_Lr{�n�|8Ԋ0��mີo��HF���b����tU�c�;�]]]ͧ������yxṽֽ�y0*�	� ������Br3no�?h ���\�F�M0��<R	nƉ3:��ׯ�9�����?uu�U��x(��'e�:qluy�����L�1w2״��#���:cH�M�Mu�f2�J&N����'�?CCӬ�����oJd�l�ߏ�:��Ҳ�6
x�ʪ�<앐����PA���|�>��
�'��������4��+��Q�%��2��䟑3lHPP� �!����.H�U�S| �9&�
p�Kʩŗ������"�v�k,SM���HJNV�"tW���/]��t��Xi���,f�W܅ >�d@�l��+#�%�y����*��jǻ��)��/)���b�US�Q�q3N�)��$�qU�;��9в��^�uO���ɭP�%�(�Ձ)r�5c�#%�uK�6�D���)��"W�K�Јw��D�ZYm_��)��>���/�.�(k=�h�h�;��nʔ*�{�k!S�l
��.467�\�ARݠ����N,edxq~Ho�/6�DNMM-B��6'#O�E!��6���:�JF�w�W�2������qQ��ߵQdf�1}%�������{�OLkW�z��+\����M亼�� ֳb;e7i����&��b"v�yb�1<�RgǅA����L�x<�%+�pUf�,
�h��Q��T�B's]ȇξ.r^o��v~�i���2w���Ԏ6+o,Z-��>[Y��5��:xd�:�s���|�æLP:��$5��'�<'ڔ�m��1����X��k�A;.���:��NRy��/��YO~9-��&d{T�_L]�ۗ��B=�~����79�ˡ$FQᳮ���g�Y��ٯ�0��K��{Z"�"E� �=[܇��9�1���~#���tt�������u��b@��<��t��-��6�
PD��C+�e��d7S�OT�}��rRTh�_c���{e8���v��@�W"ܱ�@��[�OU��$�I��������BV^�r@�&���+�r>r7]P��QӁHx\�*��E����F�ƥ-@�!�(�K*':y����GF'�[�{���en�K
n���?AE���z���(��|���[�S:	(ȵ��s �:[9����NW!����8�FK$��]���o]���:���T�??_=�������(���\�0W�K�N�
�-qa������1���� ������h� ��}�8I���t�솮�L�kC�|xě��L�%u�G*���;0�� s�b����#a��q1�۵�ȶ;�,q�ͬ{�V�uڢ;�X�T['tU�9@���0�U�z9e�re�ln��(��	�֣�P�>@���_���i|C6b��B0��@
U1SK,|�y��7䚔�`��}�����u��_W�{{��;;;��r�;�T��y�y9����V������S^�1*�h`x�'�s������p:��a��Ȝw{��Rߍ�p�܉ƂΟ|@d'~�fo�,�`3�_d�|t�KDҘ�N�k�i����'���\�����ǡf��7u�G6f�Bi��SƓ�y^�I���Dҥ1s���g2��IM1��:���'u���\��ӛ=�πa���܉��jE�<���m�.��K����EQhD��J�����8��U�o~�f�o��K�s}�>�gP>�X���G6.����S|�?=�SpO�4���.����PE��,t��ތ�@�.�إ � G�?�`���8Z�^&E�.ʀ@�\�(B}� ���O�~�Y*7�	X�W����ه�g�ϔ�����䉱�ވS�7����|n�|�K�9��������3 	M�����C�;�J�ZNˢ�`⫘!*G��^^���݀�� '��ju���Ս�����]��������yz��?J���M�M6ߋ�>XA��t��u+PχSuv���?����^����3߂�x�tY����m�ɫ5M�/gP����8R�(�Fq�����}ȷ�.�<v��۽���-o.��h�|�[�ĥ�a�98L����G��y_{���夛�$��ew>�X��щ���F&S�'5#U�v9�������yGi�|�G�xy2ٍÆ�b�/�n']�s`��ۗ�;��Q�/����.��/v���r<�	�
���������������f��͉}���&%���Y>uI�|�hC>T8.��^�,����{��V��^�dk�N����uz��R��9U�$�j������Hv����F��/�9
U���ӥ�w��X�6��7
��p7�շEo��[�`�8o��n��1蠳�k��4�/��S��Q(��MB|;G2Q0�*((K�T�Pۢ+����,4�
aLj� y����ڒ~W9/a]J������
�zx4}s������k;[[ǐ�R�v�Da��i�92��(����;x�6P��2�7�J��L���k?�d��k�W~��J�礜!��(Xw�9R���zk���wUu�`�o�a���]���d�?����A���3pY'���?O{�aC��ޣ�j��"��h��;OOOWO�tø.u�aVtA�u�>��
"�?�?�J �z�W[W�@���o����k�Ú	�ڷsh��*؋��C���=))���NZ���~4z�w�������Ӻ�Zё���D-�o`�'Rd�Xm�,�����F?��(���� ��0���Z_�a��hn��;z��A�p3!6HT̥�d8��m�kӻg۫JF-(#[\�dJ�L�d�e��*%4qP���j�n���r���8��o$��5��`͓����O�1��$֏տ"S(��Lu�����z�O������=��҂ba��nWť#I�Hb�{�'�����)�D��hۼ6���1�j��P��z����ؼ�z�/ج=���ǱW0�*Z`d'���8m�������R�����W��t��^3E�ɾ�K��aqN�$��^���즲}#Z0�ڒ�8*�6(+%,����G*C�q2~��N��%,�'�	��68�F�)EP���<����@��?.Ve�b��=J�� sx/aA�r��D�ެ�+
�t���Hf<$:ю�Ѩ�D	@Ǻ���c�Ji�ؔ�ʽ�*L�:�N��o�DOžڥ�$h^Tk����"�E,�s��({����������s"�����Or$%N[}�g�^�L�|��
�|��Ƶ�>���>���P���]npR��#�Ĺ��Vh/�E��m�+9�^�������ሠP���9�P����.1w�	����ǃ���������^��N .����
�:�T?�n.;�Bn��|�*�����<c��Xu�ڌ,r��3E�=yW`�I��E���F?���s�$�X����2��I�'ԗ�0�do��0��F�峦��K��k���}+q�� �N�&�'/��;���f"�]JV_�3��vSw7&���*��-�]���T޳[��\����D���,���q��H��(
��cL=���Htl��=�ĶK���eA	j<�s���9As�gx�v�]\NW����w���w���)��c@�v{&9�8�h�ݏ�S6T�{�п��>99�T��?�u�%������(��d*@�x���nT����Z�LM{�<�$��"]�c��� ��y�n�7x�ܩ^K�g_��Ӫ>�{O����JZb)7��Y	>�6��^��.W�l{���eރ<333RRR�忦�9�`&���9I6�,9�m{72��Zw��w%�ru�Uɠ*���`�_�D����ʸ��ma��@�y���p�J���,ߑF�\	�.Y��g*@���U4�O�l����gi�?�{��E�2�Z@����󽔡�e.Ϧ�y����iw�P
A��<�oZ����,�BVDT���x�j��&2�毰��:#|{�VMA`y���(��J����f?��@�<5YCr��N���!�W2+H8כ� �,	�_oҝp�U-�A�O��wc�3O	���R�����--��y6�ˁ���bL��L���D�k���9�������������nM9B�j�@;|ND�ѷ���R��+� ��c�3�VBx��S�RI�	�l�����Z�\�lX"j���I�9��=��]��_�,�P����WM"r�'_�D/	B�b]B6l�ݣ&��&���(����>�S�h���L���BB�gy�Q��D`�C�s���p��-��RG�\LG��p:t�U�����°�;a��!JF9/���w��1�4��ά1l����	vڪ?�3?�(�yİnh�{S�q���Td�/>�Ytˁ@�g����X����K���?��a���Y_-wv���$�n&�n�1���׿ݿ.,:^LJ����%�Q�0��r�����������>�^���-N�=�=[�fɢ-��N����K��.?%��F���%n�\��������0�_5�?��V���
fHSs�ş����U����� xq�=]ehx�����.] ���D�J�����=T���X�U^�����$���k��㥭������	l���_�=��	���!�lռ��T��V���iUa�����x�h����Pj�8^�����Fw{��|g-`c�����{٫���j�g�����'��������`������?�d���+�N�£����盛��w���L/��Q$ށ�\V�����/J7�j��<S�������&Yi{���\��CQ���ȑf�$�f]ҕ�����H4�V�zy�`�����;[c4��:w�˗:c�&��n����R"^�.�M9 =o�
�22.r?��9�bd�q��>�%���{�6�?�� EX�W��������rD�xM����a�C�)S��ُ۽��}1�K��TTIT���@	j��]�Ja���;-�Z��]�ݫf�]�㋿�竿�FC��߸��턅�����o
�����@�J?:����KZ�az��~�P�����e~d*�w��qFB�Ym��M}����%�D�JLD�5g7���4�?��~�A��6���3 �k��4e� +Ύo�U�1�OX�eo�۾G$��o��!��JSP��'=�dLd+x)I���{lvy��N{��Ј|�s�ӑ�h����(@���Nwj:��sP��[���L����6�{��7�+����j�%�m��ܩ����O0���7�u��>';�鳹�y�"=���	�>�:�&����w{E͡p�}���xS����V&wv戻ZYY1k}_[S��6�vΕsI+�� n�
#=��8��F��I�������-(�����f46��Eb�M6�U^C�t��:.� �W�Q��SV����{�*7Z�)n���d�tѭ�UP�=ז��k��2���k��նH�jC���<vv19v����I
ůU'W��F���|�H}Z�3�^�5A�!g�<L�'q<���e����;��'������q��້HnٖV��A)�Ut{�z�6�+��*1�;?_э+9@�.�p�.ܡ%.�(���ߓ�&�9����deo�Pn���<YZ��vZ��aX1�XDh��N_���A�����Âqxh-{7�璗g���%�蒻>�U�*�]]�=�R>k=��I�v32ٲӿ%̛�rppP�Piiq�G�^ � ���2�O��C�z�������� �0V���M�i�ɟL�"}�t{K`��V��*�a��m����d�K�&�H�]�D�`ܱW�a��4��̖�--g}��ŵy���0L�������gܴ?��^[|��J�S���Xo��ۘ(���G�D�{,�5��X����9?�x�fC��ړ�F�&�ع�a�����^4���� k�7oo�6����$X�.���^z�I��I��O�r�I���uP.��8ʴ�उft��2Ee�3��ގw/�v|����c���C�$*���ּ���k�7��β֟��O������q��SP�s��v�)O��'GnE��k�}���2鉟>�Qnb)o-ת�j�?���Xp��vF2�v6F�y��~Z��2��T<	q��O�h��(
���&���ܜ�B�_(D-wq&����e��h|2�d`,��?�12�ss>L����*cQǦ9�B-�yt9@
��Z��./)�+��~3�pkd��G`��˞�G��h��9a�Z>�&�/��aTK�T�t�SY^����&u���S �s�Z�#1w�2�;	��J��]�F"n���t�fPkG?�O�}�}�q�a���c�1T��:G���0�c�sF(��2����
�F�i�?��^��+Y�cy�c���:� �qG�M@���s�!�S4��rn�g����/�V�#@d��]4;;���]��m��!��t}���il#�q@�c��V�Z�[�������xfQ2p���i���%��F̕�U��ձ���e�ġ�p{na�@�������S���C[A.[d�>`zd���N�p����}�Ie+��ҿ٪���+���k,7w�R�8*��%�FR��̾O�"�c��ˇO�{g�B6/ꉡ#��^�15�ʂ�(t�c!9R�N6�����c��D
�9zF�Pj�����/����&֐�a������ea��qb�������[�F��B�a�%lLLb��l� ap��9m+=^r��g�p_���N�#�9�E=�YFNyy��E��jG�^�հ��t��UUz�ey�f���s�r9�B�Ss*��Ɂ���;���Dj6P�FE8��e��o�@oo�c�����zX��� _Luo��&t��������F�����l�^�1���z�4�v���Ӽ�r�.	���'�����(^�h��.aC/E�{�E���~�ҫ�+�B$w=X$4t�0_��7�.㝪������b�0�����͑V��g>= �yJ,����f��\� �
�Y3m�,�+�۽�XԆ�������6���*Z_RNV����W�Ʀ&|P�mN�f�Y�i�-.Wph'��LW�N�t�w���lm�s&��k�a�&ç�SE�W���B���ݾ{o��b�9���WE�vwwCqWE������-��M���a�}���0��?̤���s?��e��ԋuB5�0w3��!�=�lN�"j`��^��#�3v��_؛HR�ԅiac>���aD����!����V�9��R��V�fX'~a\�M���9�+N�U��D��ꮉa�À̋p�ߍiILq���&e�U�]����q7ذ����8���i�"%������؊F��O(>E���:�tu�53���>�J��*����&|�TI芎O�߹B ���x�2�=f:�Y�5L\o2E��3�8�:/�Ud�7��7�.IET޳�}8"�)��=n� y�j����ߦIeA�1#�N��U�����E2���QE9
��σ��Y�T���g�������I��?�0��+�xF&t��lHl�
�{��U�읠 ����k,�$�~��8��QK���Y�$�UB?#+�VL��ǁ�M�RjMН�w���ݙ� -��� qZ�>+S�)	���$]������cun�j�#�r�v4(����4� 	_�m�6��ۉ{$ŕ<Qo�
��5�$�+]�b��q�̢��C�;��(M/-oG���1�s�(��}Ό�	��4����r�������ĐJ:��J啙e�	�eIg��wzTZ��M%��B�5�{M%�G�l�O�˵+�Z�SpZ�
أ�KS���c�h=�v��ųG����ǥ�TV����E�#+�؟�����$�vS�r��O�&��~$67��HUay"ٍ�FѺs�m�4��~҆��C�1��dt	�\��v�EY�e�Kv=!���暊����S����R{��3bʈ>�J[���W��R��<��P�`>��ڒ^
��hz�<))�)((TC�<�y��V�3!�FT�s��5�-�(Ux�"4��_�B�>�$VI�^G*�n�bn6�ü���dG��Z�H!P"O���7�π2����CG_t���s��o�LH�Ό�:=v�/�Z1�'����f��Wf����;�8�� ����B�G���6�es���m���궘�n4��
u��Ȗ���Pq���E`o������4֪@���1sԣU��]�?�n���~?"*d�H�z�{�!6�?��8��h򨉆�D}#�4C]]=����M$�V;���7z�ѭ�_� �HI?�q�].]�/qpr�]Z%TS؛>����j���;��_���,}X9�<8��*�����R}>�=����Ġ��:::��}mĨA��ɡccԜ�
�og�X���=X� {*E�=m��٘e�Oso��c�Қ�Htp�2�����F��n��u�������NC0]N�F��=?Ԭ_9�=m �x��ch�  P��6o�ϋ�B:�[�I�����������]`E�Lϯ�G��>&ڵ�X�����[����
��]̨2��Ue�Z�\Q3An��3y�h���������Z|�Ȃ�B���m���qpRl�Td/�l�oB���?{������<�,�4��k��2��:=M�V�>��|>�>���xtaM4Wo}�杺�!�Q'�{G������
�e���1����+!O�ZfSeb����2��\"����չ��x�%��ٌ$��0��fӌ,4�S���3�U�Q|*�	�O	ڬ���=f�f��?�cՉ�/:s�2<)��а�7�u�3Q����̟���y�����̌�
g������|�,�d����|ڰp�ٖk��㜹�s���\��7��Z� �Fٯe�^4����o��{��j��V+D�f�5`�`f���,m;14��D��Z����E����<=�Ҧ��!����+�J�'�u��u������bؙ+� hbcc��y���>���� ��;�ey��(a���7L�8!��r|��Y�Z�
@��0�[���/%)�4����яi�ҏ �!�+�saʷj)'^��"|���R%�B���eE@CI���w�	"����_+	� 2ݲ���sU�Y%7�&V
e��܍�*��'�-���XW3͎�/���b�jiI@�����6�0�~���U6{���i{���̈l��OP1�`/��Ƴ�z�!s^^b��hmt����v�D��7E�M1o	��'��-;�v���P��gS�{Du6�;���_��;�3g3����V�ݼ0�ۿma��9���(�F����m�5���[2���S�d���{��[\V� ���V�6��0�]���� ��� ���@^�d�j�,�gi��C7��1�H	�S&�U��o.�(C+)�;�M�p�{�_1�i�֨;5E��+bf�?��N��h#�6;�q��#JdP��<G&�H��=)���$��g�"-�E@rƕD�P��D��j�Y���"d��А%��@�D
�������s���TR%"��"�V�[�y�B�b"�oתnZ\���"4��7�i�y�����(]O&�;��z��'�}���E�W4i��೓���B�
bM�2�?dKj��k�C�Vp�d�D@�m-t$)��RU߈�'�c|_�q�3�0��	l�9�����>��ҟ����s���D��ھT�#[�v'B�7Y|�c@�`��s��ŧ�(���" �=�id�FgIb���U<��Y�`��h�?W�Y"��닇%� ��Blo�3�B����p)�&vr�����ta�������;�x���ܩ��
}�oh8ėڿ=��HRU}W�[�Z�����$��wi�_���\��	j�t�@\aH�ͥ��}��'wxS�G��uiBW(h�,�a���}͐*h��V����P��+O�
���I:f3N�e"ʀ`�!�

�,&B�@ࣸ`��ה{M���~Y"@Q���5��>1�:l��M_�0��^�×P��,_k�~��,�*eND�&!5�? "d������+�qP~e���w	;+���O���~}����~r�2��Bl������ev$�q>u���qq^3��\O����AP��p����PU�vL7�� ~+�������](��v�ቂ�1���բ�p�۷I�g�J��Ƭ����߿�f�v/�)|��!}����n!y�Zᩬ������WԔ%�=h�[���&'��N���H(�*�d3��N�!�Ƭ�O[����[��,)p[Y�$���+/j`4�W�<~�����C�̰����>u�N�?�H��� �d�`""���B�%�k��˶�>�Q����\�`ͨ�Q��;��S�K�g�����x�ml��"�Z�^��J�"�A��+}}}�7�ƺ�
ִ?�l7R��3&�No��NzZ�@]j{��ϱ=-�h{	�%h�s_����L)�0������-�{G]�2V���Sz�v%�(�o��f���,D����C;JDF�\/�,o�Z�u-޳���~2�
j��˸��l���;n�qMW�K�cF0�Qi:�y�ԁ��@,��߿L�Ʈy*p��/�3yĳ���H�%
��y<G�x{?|I���<;����h��E{2��S�y�?&);�~�{Gh��pz�4$�E��B�e<>�������a?�g�����|dk��&��y��^��ST`MloI� �%S��vvT�o��:�)���p]�����ӣ�q3<�ٛ����~�;����Wuehr2�ޑ���Q��9�633C�Z(�*�����&'Q����Uc��)�{{C���#����������#
���e����,���&`\jC
�{�`�S` /%���aH�m���ۮ# }��ʞ�؛�+��$p�<Y.�I��e{�!�)�e��"*R����LJ���C�-�C���ݲ����7G��/��}�<��뛛}<D�TM�JYlT0�����ڟ0˱��o�*'p/Baz[�)ֳ�6��m�$4<$/?�װG�8ۉ�k����ڦ�Ąp1>1|Ɣ���jߛwh�D\�1�FO=W���?H�K$����F����U��E��`/Ow��u�$�q!��$�X�5�9&&��߬��z�A�\/j�w�T�?��N:)@w�78 Z ߜ�kM����6��o�_$���l^v��F�2=x���>��F8P$Ņss*����1*s�з�a�+����At����2���fВK�:�򟿫��jwttˍ�,�z&�OV��Z ;e|��	��[��aC�NE:MD�[
��eC^4t��A)���O�uX�; ���&���X�C���*��!"�%$P��%N��Ζ�z!���=y2��?u�4Q\�=�הwJ���|$���|#�2�B��UG�"B�?^A!(@@����V03�L��*�[�"�Q�+<���iG�اG�m+^�\�>�W��x�A�6$���5G��7>�QZ>���P5MR/���n�`��q+J�+�/�U��Qss��Cv�H�n�fH_���U;3]e�cn	��[U>];��//W�?5%,�41��E�Ã0�-�*�����b����e���eHeE�4�Qu#.B�ʚ���l��P��~�g�V�]�S��k�Ơ�Za���A�a�p{��]�#/�5�?��aD�o� B+���pf�QP�J��T2"Q.n�#���%k�N[�g-����Ȁ���ddZy��7'�y�݊�u���?t���� �S�%��û����M��_!|i<�K��.���C�����m~�?w�|m�7"b+��o�@�Cv�c�`���l�!���A�+ �c�s./l���yQ~aqi�Hb�����<aaXEڛ�Q|��o�j��`����s�{�v�(���ʃ�:��� ��-fc�ȄA1��N��~�/1G6k?-/Ti�j>>T�<m���/���ݛ������c�.��kk�v�ެx�Q��?�k��b�SBQ�*ʝ�s0� 9��5w
f���"�Q�pRNZ���3���ay��΋#��a��|�2RB�U.���	/��_��p��3�Z��>#I�&���v����Oh����	`  *2�Z�94�b�WDzz�-絓�S�@tU/�� �ܳ̓M<w���?��{V�63u���1��� ���0'�f/AGȥ�����P@NѶ���ˍ:l�F&)��b�����V�m%Ԗ�%(@�}CɳEW���9t��n�O�/"˄Q�`�H)��$��P� �������\ct��������d_Q0�7y�	Ǖ���t���2��~���M���{��#�gS������5x	��"��'{�l@K�@����%B/ָ�&1�l�=9������2��d>�W9��%r��u$r'>�Ɓ�I>!HmDvT�����t��O)�1�IZt}���2�yklys#�{���hS�',���B�S
���n8�q3{(�Ņ��2�Ͳ+4�t;�t�� =�|}Ǎ俪�A4/���
]�\��l����g���p9�������hutr�0V���K��*��/�M];�����F�CӼ����V��2_���qQ�%�戁I�W,+w�W�����/H�+-	\�������M�_PR 9��O��yt�[=(b�{J��ʘl�R�~������/��NE;��a���*����ϙ����A���H�|:+u��#�O�f�+�3����`�P��bWW͏��	w?��� ����Q����sUP�肬�@�����ME
��mͪ᪦o�Co�w�a7H\�Ba0�jIIt�����k�Έ�A�-W�}u���n�RmZ�;B��5R�/����r��������xf�8\J������"�j"K��qsy��juә���^\�{��;���<�n���� 	��ҥC���.^e%�G�d��P��U�ty[�#��~25[������j�g����Yff��
�����8���j�H~�P�!6m�������2�6tKn�A��1
<��yoMge�KiQ�R>�eԪ��o������L����⡓g`��YA���烩����Z!K�O��$D��RW�ķ�%q3����'�;l���0�u�_|{���h���/&yff ���Q�^��[�;4aтUΎ~�K�������a����t�����Ŷ�Qu�yq�eV^m�hPP2�R����Gje��1��~������!wk{��Db�$�ɻr�Z���V-���?���eb��m	yޏ����8������K5��͡*�>D�,�¯�]`-�K��/��^Y㌵ˁ���i+�Q��]�\� �@�Nƅ�N�;�2�W������]�->Q�N�����?�x�Oy�������ο[!}� �+�+*kmJ)in������'�D�f]��S dߤ(,ܯ'�ⱙb	J���C{Ǜ���*o���F�x�a�V�#�;&�j��7������	A�1�ū"[��E��h�^l�ƕ��m̶�3�J(�Ύ�F�r|bk�����WEݙO�Z-~,�.�
m<�^���Mfd�?�{g��$qL~�����L��k#�by?w��(J��������`�}��d��(���(�x!�e����C�$�9U17�
sht�x��>ݤ���lg�߅��7����R� �?3�:j*����Ƹ*U󺚺EX����yz�,�x@zI��� �@]���{r� �����y���޹swmmr|ȓ��wڶ���������j��o~���t������K�<<�ήn2�ف�
?��Y��J��；�4� �<��
�"�+ �� KT$$���#�I	@��:!���$� � T��(  ʠG Y�A�E�Zxph,k4 �	w=(�p*��T �)��+ �!E��lT�h��(��ιzQ�^�MO�un�j��������a&�!������|�h�VXn!J�)۶u��&�9W��9W�����˗�O������h4�|yo}}���P~���[�[D�{~X���|~�ڵ���[7o^�v����U�4v�ιh��<6M;}~�v�G?�������7���S�(��m�jt��Ս��(tmw�֭+W�M&���ѓw ��½k����>���O>E1�Eۺi�)W #+�7�4
^����<��_	 Rj��ʫ��
$����''V�#�KХ�B ��u]�}jޑ�J���j�.#�!�o�9�w74\\�7]�|������;gocŃFDs �f֊ 9A��3�H�u*��}�Gfi�VDPbr�Ș]6�.%��j�6�uS7mk�:bdD+񑇏=�,�9��������g�������͛7����,�b{k������Թ��~ss�޽{�.���ի���勗�����fU�D��FeQxK��r���i����Yi�B���	H��r� ���2M���WªGh�{% �`s�Ɩ������.K")��T;N�)�JG|�b3o:Et�#������m���[��d'!5�&�D�D�����T�h6�-�ES7������v}���o7n޼re��'� :@P=<>:::*�뺮�{I��h^Jz�7MS䡆�eŉ��K�<r��e�Lr�d�%䎖fo�z�43�Q�w��*��Ñ�6���*E�pӵ�-�����*��Z1 8r�;U�A��*F������}OD�b=�ҳ*0+�Փ���Б��=w�,�4T{!�r�d����!�]-!b��:���J{\]�K���xP�)"��:"@l�nQ����$��+aSr#���
�]מ��<}����T�INNN������u^�?8P����'�^�zy������ͭ��ӓ�!R[7P�Ս�7��vwv���q=_L��v6w᝻�lnn�|�Q�^��ͷ�e����{�̓����V ^�\�mU�ϴ�y΀���Ƚ#� �b)c���L���~�6��n��f(o�*("�gn:	H�=:��h�?��"��E&�O��L�z.���鐭KvM�ɡ+J�*JV�$h�{`5�<R�PR�!}j2[C=���Qv�?83�M���v.q�Q5�L&6~�{ �*NaV`�\UU�ܵ��]�F#�h�3��)��������˗/#�>vO�>�Mg7n����D�Ǐ?�������NUUm�UeE@�ɤ뺃��2w߹syoo>��]�B�Ǹ�6y����ܾ���Ӫ�LKߑ���˪a�����d<��ڵ�����W��y��W��y���b:����z�j�����nB(�ik�2�OYegg{m}�y߫��ŝK�>���Ǐ��e(|`� "��ykЕg6�w�b���'����?�J��
����)���̒�Y9r��0�cOE�0 �SH=)WX
�(��巾��
*����'�\�s�,�[yv<.��o�{_��Qo��o��>�'#��u�ȋ�b6�mmV�5��1F�<Gf������0-U1�K�۶������w �"�@HA���!��:gm X__�����A]׋z���#�{ύF�w߽KDO�={����lZV��tm{��O�&}߿~��Ν;D����E=/B ¤h���2�29��.����Z��R8�0!d��Ys��&�L�,U��j�����B�|��x�x�,���9 X���1G*�p���l���:�<����CTD�!U�;G��1:��Oe+"�9�����Ã�T������+Ua�kk�0������{im2YL�����l9a:�,%M����\0x:(Z��%��T����d�gJ
��H��,��0A9R�._D���y1���8����"���bQDT����'��s��#�bk�6��`uKJ��5ȏ�ioQ�����1�؋R��w��}Ep�2��
@d��e�� �y(�OgW������dsg�%oֻ)����6}�-G�d��ANJ��s�,�hT��;3�T@jb�9�DDD�����|�P]8�����˗���[Uu?��7k��.���{��O?������?�w�^���G������k���흍����D\__?9<~����K�/�^�u�v�nomM���g�Q�Q5z�j>o R���j�8g���3���Bp���L̤�b$r�����̦�ͤZ+��U=�Âֶv��3�ͦ�l~em}��
ߡ[0�^�몀��"x Pa�ʁ�>�� QG����"��:1&:Nb2�\9$�R��b� �e+h2Y�\K��@��-ꔊ�T4j\&�@͏1�s4Ec�Φ]�zrλ>�9{��VP��e%l"��99=i��{$t������!����O����^[_?<<x��z6��U9�M봪���k�0�ϛ���HD�p2�"���UeX,�MY"������5D�z��dmm:�����@�DD@��18x������g�Ν;���7/�&�(�z�~��������{^[_C����Ţ��PaT��x:}}��{w��uU98<�����������ݻ�L&���^.s� �y5q��T�%	���V�J�`��S���5�TE�v��/�����"��������:k� lI@�φ�Pe�K��OK�jһͦU�A�R�<�eSDB\��osV�w�Z}`fU���w{Dg�̜j�X��Y��U9b�#'�A)��,�0 0a"V�jlsP��w}_�E(
k�4��W������7��qJU�?8(��4���FY�GGGO?~����Z�9�B5O��'��_�M���+"x��q�u� �*�ju����Na��#���d��Q�#�F� �4 �杋*��"�Y͆�R���H�5�#�*�1��ZbbE}���f��	�k0%Sm�#̴���,����VE�QUE�/^�2��x<^�J0�e�&�#�����yo���'+@
�ڷ]�#T�C/sY���ŋ�/��TЗ/_={�tm�VV�xm��ʮm��#aV a���X�&&���C�\P%�pU� �����yR�P�s�HmۘB0-X"TPG�
b�:]�SZ�+��9�(�B�������8r�7��n��!Gc�]j�K����ܧ�1㭞 #!(p�D���A�HuJ .�Gª��,�嘍vn���VS<���P�DP�5}�!ϥ`�M`�6� |Q���!*�ďC����&-�������l6�뺮�뫪bN����˿�˿|�;���M������,�O�>y�4����hT��ӓ�����ӧ}�_ݻ���ظs���˗�z�u.��o��y��m���g?�r�ʿ��)-�glk#�R:���w�rM[4��U+�B�4	c�  
Q��T�s��Ξ��>X�Nw˵�x������g�����Z(��Y;�ԱW��5�kۛ�kk�qcݷ��ʽ@�Wn�6P� �r����
�J�$����$Gj����)=�x ��*�* K=��܂���ʑ)��SՌ�*!EQ��c@��;�A�Y����TWD������׋NOO�,�����%"v]�����^�ƣ��ONNNq:�/�w��lk{�i��|^׵����?}��{~p��흝����Ǐ=y����x���f�Ǟ��ݻ7O������A��"̌OV&�L������ȹ�g��֭[/^<#�Ѩn�y��Of;����G����w�����l>[�\�����\���o?~�s�R9�^�z5O��7߽���~���K�[�;��/~��:�����%��ت����Ċ?g��+��K̀���y�mu�d��W�����L?UBZ=J��"�P��������+!�o����g������.�k�R
,
�.U|���s? �����Bc5Ur�z��)$t�ڶ��������7�O���WU��-���+F�N�ym�f:�.�EY��]�
E�9�*i*�pDIt�nU���Ǐ���;���Y]/��������Y��O�S�����L�(o:b''�6�!U`"\�!�����ʋ��ό��4yI/		�p�,LÒ_m�W�	�r9�hzS�H�-�♭N��9��PU�e( DPc�Q�R���ah�d��������!!E�v��=J�> BZ�6i�C���})�@�!��>�M��3��2�	�P��ٳ��������������n._�����Ƚ|���:�&ʇ���J�|�%��"�z���w�0FVU�<�+
��r ����Ҩz�M��m�Ѩ��Q�5�k��h��a�d�lCeQ�P��%�ީj���<��euW��m�-�. �Xm�@r�2D�'uD���}d����5���x�iN��`f�4kR�Y�`B���NN���X� �ּ<W���w
9�]c��������E�L�C$��xckk^���������P�~K�����Sf@c��W���%
�(B�u�E��fY������F�?�쳇�m3��h:�F����Ƀ߾|��$@@IA�Yu�<�/��H�1:��sc��TzXe�K�*�ޅ�d�B��� "�w�ù�༖�V�QSq|�cJ��&@E$H����i#�S�M��i�NO�N�k�jwc��p�=��'��/<�pdEVU1�h��mFD�Y}�q�@J��r�%
9��3g ��,�9���}��M�6]�E�(,"�#!)�#r@�s C� s"���}$g���$Q%��mM=��,a�K���y/��9��׿��b� ��bqzzڶ����#�����ٳ�|����\U�#s UUݿ���̦S�Vɹ|ҧ��*�0�67��o~�������?�Ϟ>},,��|�siw}}c4��h�t�h��w�xz\�MT޽r�����-�|��G��>><:�ۻ:;9���ǣ�O~��~���?��� `Z"IX`p��]+t�B- W�*(BJ^#�vҶ�S�巓���X;�%au�9���RPD!��W]����8�ʑ1�<�!&D z�P����tgg��6+�_�_��<���^��os�R��g���#�����EY�U�"�c���y����t�#QI̳D; ���ɤmQ�E(�REY8x_����3a��5�U�{O��u}zz�NS�y���"�_�ΈB�bMm�:�wC*LR^��3ѿ��p�_R��޽:���������
t��uj
���;���̺�!"%�����i��yZ�H���o�q˿!��U|� �ݚG���Rvqu��C��D4Y[�F�baԚ�(�śt�y[�p�&�0�>�uS���(
s75E�Y�5-Z�v+��d����X,���["���TE��|6S Dh�v<�h9�i�d��iO�PD f��0��@ U)RUZ����	X�*gf�}UUm�b�ұ�c�6���7D y9����Bp>K����j���Y.؋ֻ�(/1d�K��-"������ |����9���	SBm ���}9�~��d�=�Lp?����e�4M��'D�>Ʀm��ca�)2G�Y֬�	���ھ�u=�/v�8���gr~�t֯25P��n� ��"a=_������˿��>�صmӴ/_�l�9��m{z:��f��VDy4�~�Om�� ��簲�Ð�N�����j�pLT"�Dv�I��W-z���ӃW:��XlW��j<F��Ɠ��iT�w���9���F�t�	�Z����fgg[�ճgW�~�Xt�4F�g�A>��[O�����R���_�X�A�թR����<*Kl8D�j�Vb˽��lx&h��l��aLf�	�����|��]�aTUHʪ(��d�V%3H8�Mì�}���QQ�Q5�M�am�
�DސV
��YU���d�������iQƞ��>z��IB���Ţm"g�>!xBj�v6����T0h �-f���!�w�fӿ��_��������/�������>^����+r�����~<W�����f9����.���_��/�����G�|��xm""����o��}��ݫ�/����������,/�oXPH:o{���N��1���AA�v��|�{{�GGG��TW(��L��)�2&%  ��� 
�������.��$Ul���(�Z�;�K�2���g��
�1?텟�:Ԟ�\6/~6[7o�@UEL�;�~�Br�9��	>�1��Y�j��LSPV�;g%�&�j��N@a�c�CDO�Y���a��Z��]L�T��z�l�"�).����3�+K.r��cF=�a��V���5$�1q�T$��s�h(:��'��%ys��+޸�?g��d�N
�K�� p&�s��!�Q�9UU��jU��s���)�Taj�� �v�+@�u�2�ʼ�/�ә�+.Q�4�>'!;�Q��
�Iܑc�U���XH�juUZR�˲�y���w�:��t��q6�q���|[U�[��y��&�B�����fj��0Jc��d`25���AAY�H�����։y��VN�4�Bܸ���C2��7 X�\P�<�ɳ�W�G�}L�;�Xm�r a��* !y��_SpFv��`i��W������mu���4�g`��'��޺�V�8r ��}��>����*�	��:@�� &דE��J�K��6�Z���j�0�g.�D�E1�FmՍ�ck�鈚���){^W�u���u����k}c��~90����9�� ��3�� ���]�]Y�� FZ���4nSSl@R�[����	�l1�������W���k��M�w�����j�<b��y���4JU�eUqU����M�0循�+ׯ7�y������ޞ�'���n49��_?{�����Drs_���/H��ק�fZ7�GJW&����%˜4,�z�Q<�s���=F*V@B�,�J�aō@ľ��,KDUU��Y]+�x<*�����-�/}��
��@�i��6m]�]�Ef1]*�#BjaOd�5������|>_�MZ잇8��������##X��U  (�!��e��d汲~�����������������k��������ݢ��ܸ���Q�������/���w����_}�h���T��pxp�W���U�Z�y�ҦBaB��ڟ��f��5���f���/�,��y�-��9��c+�]�?����Y��8F����l�^�
�=�#h�c�u�ୀ�C���l?������������l�y�+��_Ò2�F���(��\m(�
�""*0�y�������=�)���Xb���,D�R�q��h>8QU��u�B!��h<�Y���"�Ds�[�$he��	mKe�a��:e��]�A��YZ"r����.[y��2G ��(�|8�X�e"r�] �/V8k�#�}4� �(f�1W�2�('5��žE`��2�$�@٭��`+�E"pn~�pz��y�I�)}�e,XS��ÕZj"�0Ї@����~mm�t4��\vH횓��*��y ��&D}<:2�uˇΘ nnl���x�wv.�h�v�[[}�#����{�����믿���Ob�`���xvԍІ�d$% T�	W @$PSk5E���9��g��d�$���ZC�Y:6�" :^	bt��'��(ml���
��r��c/�bIp�st%(JO��`*�+�ɀuM�+��@ Gd�8�* Y�Ú���Kn��-��E��Ό���SS2�A� �� �:R'p����Ͱj��:��r����@���<P
���;?����w�l6���ֿ���h>�[���^�6���}$$=,C�%@B���e)�tZ�:'
��ɱ�_���j(jc�T����	�J��
dؕ"@4_)
���
��ly�xg�֨���W��ho<�@q*�q��VQU�6�(����iQ�"h�� "ĺ]8g�mll�e�ng1Ve�V.��yy7�;z5_4�W���uY��oc��Ӛ���Yծ F���U�:���9���D�\�����f�(����;JT����Y�Lr���Y����Ύ��ʢ k��	n�Ah�*H�1E���(󐬅�2���>d�2�<H4� ���7&h��lw��@x����b������{'��ED��w�i����Ӈ�>�������+/_<����NO����;��n�~�j\V���� ��R�/Mj �K%%4�����O��4����uyWA�0�Z�̆�߇a�����M���B B
�{�c�'Cd&B�Ot�1�06w�"��>��$�*o�) �sh�Z@6<�����oh�����%� Cܓ��V+���OV�l~������ߢt}�,�71F��yg.d���Қ���s���r�4'''��4J�V���7+	\x��}�ri�&���P��Ϗ)Cv�0���9\��L�A<�$.��+͓���V��"�ƨI���P""!�b��]N�(���D]�Q�S�Hd��� ��4k[Q��:督�;M`"��g����8o�>0������y�Ĩ����9�>��l�
�Ժh>�3m�Yɲ-f=�.���,�W ��۱�ȹ�]׵M�X	/s���!�c�-c���[��	�1�����m&�s��d���c�9�;�"�!Q-�HD�.lc��eU`����3����� !"s�ҩ s�5N%:���hb�.�Z@=����a�&9��������5�*�E�3m-EP����~�&]q�8P@�eT����S!s]�ՙ�%SA;r@�E��jx9A���H����C,i��B
(���SY�VuXU�q2��蝳�G��F�BE��pvPE�
� ������AS�jg3"ǋ��l�����*���3_U	TK�	�IY�EARTT-
��b��H�P� �,����om�*i{e����A�u�';���֛�6�4�ӗ/��bۅ�[;#�����O�<[t�����[�!F X7mӳ+'�\k �w<S���- ���tm���p�X�JQ#����d�r���%h^	@�&w�������{OHVc������!��^�5�I+ǂ��뛦���kۺi�����a(j��j���NDK��*'��	ӧl�U�0�,�D�՘sp��FD�v��t]�/�b2�"��������ϟ���O���[�b���f�kg�9+�m=�O�g'M����׏>P����?��;�x�����?t��sg#�t�[Մ���4�'�2���wޑ3tO�P���M�A3��t�J.�C��;��iM�9�j�K��������J.��q��rC..���������#�HV�)+���8�V�xy2��IZf9�$�)^�"��h�W�d�{TQS<U�`�Q�zPQa��@�w�̌�,J������(���*ZT�*&�2��#7�L���-�f's�AJ眈
KR�DD����lt��g����r}��c$E�bѲ�C�3�N�#M�g��|e^jfyoe���yU5҉s&_������p��Ui6ax]�����^�>B��.x6D�3��%q3�P��ޤy����PGNAb��;��MC&����c��b׷�r��֑�����ת�,�~���~}c���ꫮ뉨��h9!�x!T��tvd@1�93��Q$�P�j�7 r������ij�1��k��fϝ L U������* "���p�1	��P �\�3@z�e�ҴA�`�2��9Gd �:�BY
J9O���]5��a��R��;���Mg>$D��Jcv�6  �
%x6�V撕���{���`!�yw��uL�L�E���g�5:�X!o��R��\�D'QS���({�V��X �R��Sa5�BD���b�Q%#d�\GR��|�\�FcNA���`/��<�"Qt�Dc�2�*��<M&Wd,(�QU�+g���Ƽk�����ڹ|}��uݫ��/^��0����-��P�=�f�µ/
D-��X��ln�ͬ���m�u�k�;,�Ø�!��HBA_��~ǵ�~�Qp��=�]�M&����F�Ge>:8��L	���2��GT�E[D%�Σ�eUnmn�G�>�k ��q)��D�����C�,C�]�ED�t�WlX��1q�'0=4U+0��G���_d�����|�u��|�R9��'E����>�����{���|���[7���'��xT��={���N�SD,�R I��3[Ϯ�Ϛ�O�*�7��>L�a8uy
jR�c����Ƚi��}>������%a(^E�������w�7�yɖ& P(����3�#$ `aJv����J!PV͌\x��`���V����R+�_�F�f�E�hJ� ���z7���7��$�0y���@ t$��%Z���#n�F8:BUEe�q��=��E; *>��e���%d���h*�7�=��z $-d��&����1�G���! X�1Q�ͽY
aXp�qn}=�2|=GBt��)[������.�nP��;X��{��喠̞L���`�k��&�X��b�h��YT�m;��OREU6a���q�$�3��-3��2��I���ESb���˗/����x<	E���NOO<x �UY���؇��O�w+���Y:;.�Z�jK�"*�"�g[bO��d��c8��,| �h����{�LƋ�(f� ""nHU��I
!��O;m)�`�����1H����;[���O�PD�M�#�  ��T¦4�r�Ϭ�4�۩h��P�|���f�uy�bRrI�6�~y2E�������(˲�!�F��󎅃��j pV��j��w�;���h4oll�}t���5����n^�y��iN2%�r�NA���
0 ����.W�r;����3�PJ�"����hL{���](J"�(b�$5$�R%��Jj�)
;TK����ܺ��O�1r *&�uQ�j�t����b3ݸ%T��mG����i��T�C�H?�x�t]��D`ޫFWƓu�!��
bpLԪv���n踠yE�Ҍ�a<g��+js��I͊1sd.��o|���Z鈊"D����w1��ł�_4��M�,�3k?��֊41hШ	:D����9��g�@L��a[����T��`����kk���M�*a��G~�����/�&�*	i��-���mSw���2�Z���'Of�S$��	��^ID�mCv�`��O��;/!fe�T��v�f��*��\sȅ� @��;�ʜ�Z~Ȳ	'+�Y�reu�/̉`�����+y��Z]��cfkW_�28��� *�\�ЭQr��L��sg�p�+4�?l�l�S��=EDt��G�����A� 0	҉u�
ɺ�Ȣ�C 9�h���d�w]UU,,)r7O��ٍ�hB�;��c�6�r�3V���E��Ð%X)�\JQ��h��j"H�2[���5J݈�����"=�<'1�t��1�R�MB��~a쭚��7�%g��p���o^�x� �d #s�%�u�~;�˲d�i6���ۻt����ק���e	
��F�;�`��L�<��޻T��+μ3O��*r||l={���k�(,��X���'ڈ�a��1%�"��Z�����g���n�YSIY�]D��6�3�Ȧi���ｹ�f��F��Dk��Fe6s�
 ��%=fQ-�«�/��P�������w̱U����*Eaa�������$1��u]���9(��г1����m4�&�&f��0��]�~h�ncd�L ��b�6���6*�|(�D�u�j�.+�u]׋M&6:ifD?ϟ��L�$6n���"\��XSU6\�#:A2|���F�D	H�1Y�6���(v0^ta�0���Eē��p�y� %aE����Z�S)G��d�g3��V7�dH��2D��HG�EB*b�s�&�8��뛀 nlm��U��W�ո��eW�ֻfW��]�ܾt{2�8�"�J��D%b�Fx��Ee��TԳK}��~^�b��&0�X,N�Oڦ]�LNON������K@��:A��ED���3�eY��d2�,jZ�+WvY�6쾥s��'��y�$ӌ�u;�l��sp.��EU�~�rm2�Q��� �jLk���w�mV�������#e�༈�]'C�̀��X��"�"��չ8s�'��𹵾���H�b��ɭ 3�6�(`*c�b4�\9{Ĭ�yT�ɚn򢭹4�9K�֯�ï;]��KY��[�'�e������g���y۰Ya�H��gǆVQ���2��2�u�9H���4D6qf���k[�����t�i>/�ѲX��E#��;L��i���P�����xG,�d��ͻ2h�^�zv����1ߝ$� t�D���]���3���J^�J�X�!z�
g؉���ȑ�Z{�X����{c)ڤi�Nj�s��wA�#�,w=���������΍���cߧ��9�7�R�H�K���&-���PD"�9� br~��wޠ��6?�AD55�C��||\���g��̗�������׌ ��Q�����E��n!��zOU�TԘ��Dk!���[�Ӧm����R	�Y~�젝�g.B�d� �#@$�(8
�r�C(��f=��#j����]�2ԩ�GM�a)4���)/�\��k/���<�%L��_e�ZEc���eAŁ�j��潛n"��ώ�;��jT!.zU!b��˫e ӿ�����):�¤hߙ�V/�❘%�/<�2g\��D�������[+�����B��E@r�Ȇ��'!�)\
`]� Ժ7(�
�z�!2��s����k GT���H#GBE�P	H�T��b���8@���<��b˕��9��]�"̦^������v}+��L�Sݘ�K���ҳeWUU}�[TZ�UY�֚b4mlllmny�s�" �j�j�Xt�i���0%���NONb��S��yԕ;�|G�I�ܝ
0@h�k[8�9��fQ��K��Q�@��"jH��뺮�s�Ο�ɟ���o�����k׮������_�x��,t�v4t߹|g�W����;�le�fC�=� ��9W��"Ǽ�I�jHES($��b�<����q'�2��3Ê��g��̛���Vq��h��v�����C�i�t�[.Z��^��Y�q卫n��a��}GP1U�j����U��-c�Z�����,�2�PUUY�����yqV�EL�2����$�~��Ӈ�jҦ���g�Y+W�w�$\~���u��	��Ч�j��\9Љ3�p��QY�㩋�0��WƑ<%#&����tZE�z��-�"����y\�G	Hc�z>���O֘Ed����^�� �����p�w,�F.2�9G��pdu�j�W8�ˌR��3��9gIH$)I2��)��>�~��������c�>�����@� C��]��]�TڛbQt�ĺg��C�=(x ��gd�~,BU�[�жq��#
s��Ԍ�n�"uH)�O��5 ������6���*�c|+����BX��Mi���*੫K�VCV�u����g� �Ҵ�9� ���
�_L99��V�����9� "AAQ%+_@*�|��($YӴ�23m���'�1�EȐ�IDš#G��Źj1G�b:M�7�"z��|pF� D�Ǵ t09nU��YSЉ�O�����#
(i�2�f}�<yDԫX=: V�|��a$�@5"���J���2�:�sT��"Qf�T�0xf� U����M�QAXb���x2�ll����}zzbQ���{g�:��7��c���(�����h�X,���n��dd������:�T�����-��g�zO �wCo@Ukz���]��t}/�4� ����w�G?�����o~󹨬��߽��b>;x��9��H�)��o^��.x�x�*��Kj� I����PP��TŞ�"���2vC�'��u�VQ�x�8�9%rnr-O�M���f�����eO�D�9g�]�S����k��ŵn�$�)����j۶�4w���d���BR#�l �b�899Y,ɚ[���RΟrL:���A����U����r�6F��+��&�2���7���a��-`�&.	�r��q���ܯSC	D\j��c�8�c��>$C��v	���ˍ�#��m{xx�*������D�`IF  �:����J-����w���s�ڕ+�I��G Q�)3nm���("�P�
�s���<�l��$%��ʰ(9��Ȑ��.�``�s·�6���7ٹ$Xf�iZ��=jy_1T4���"����On��sޏ�U%"���+�]�JM�s� ��Q��!L���q�}F��/C�"+�E�Kg�߅�$l0�J������Gt�r�kߚ���F��Y� �eB�r�%���0������-B̭jb�`�h��V�FD!���9W���Da���fN��5  :t���i��IM)�a̎�ʶ�0ŒB�5��@{�H�Y���$o���Υ�l=�w�=
�s�sO" ��v�@����v DT&�U;@��
#GAD(Q��LH��)"8MR(ʠ�D4F�:,�ʑ�ȥ��f�(�ɋH����u�[���R�oB��a2-��:\VΜ_!"����m�"���޳Ǐ������h46GߊЬ�YY4�j, E(cY���Z��m���b1�B��u�4��w5Y���T�˜cz���򩦪H� :���a ��W Ī,�U5U�g�ϟ��޹s���;㵉�x8M��,�T�pf����v�J��ᮈ�U,&�d���P5Rr�|���w�W~��|h*$M�IqYɻr�`���Ѽ�Q�j4 ��pK���5  I	��xFmC ˑ�!�2��j�pa�I!m�U^��k�A��H�����{��HB������V,��B��P���������"}3�i,q5�aL��;=���[���U�ֶ�1��[[�X/�TW>%����Ǟ �AJ�� !U��d���X���)ɩ+�K��n��o�����Q~�[;i��z��uD���c��C&�������Ι����D�i[�B�\ ?T$(�u��G���6�i>�J�5QM��)��V{�iT�	.WD��'�i���H���ѨZU8E0�'�������l0�tdHbX������R�ȑ%�r�F�#k�
�F�Dt�(I�,�C�	07ki�p��j�k�b1bbLZz�� �J�ák�!r	�r��Zڕ[�A��
���=��L�9Q~�8��S<|Tz��b(Rd�ጧ�v\�r�5��Sp�Y�����b�X,����]� G6��M��ɊT^��ҍi�cP��׬A6�"Qr]���^2�Ҹ%%�\��T8�}��~#�^E�zX��%i=`�Ӯ{�vr2���h'��`'�u=�*��'����ч �Q	!���
��!�w�Gu�$�ő��
l��<�ٟ�F�5�&[�����/I�9[6_Yu����S�$U],/_<G�c�v��&��;MG��w}7��M�Ӫ,����H�R�[�x-�?	��sѯ$\�ɡѤ���{O��"�j캺�;��ܹ��6�s��b>��u��(��&��
I{!}+`.�R'"�L&]� 	S��'�.�O�9#4B�Y'��X) �~���.���)W�(�g�M�R�,���Ȭ�����=��|� @)9�<�� "򒧅W����r�	�1�E5�ƹ������j�E��*��r_���+�m:pH �s1F�$*���f%8�� �8����Eb�f�9c�dBo+~��A��������?�|P.T���J]B��S$���X���H��4���6���2x�\�d%�?�.��F��#��O��N|�����>�������m�"}��u�4Mz�ܮϖ[L�X�nQ>!�1�>��A����3�*Y��1Oip4�L��&^��D�q�3o���q�Dn<�mYU��Y:��Ua��ew'��xH�A����A�c�L�ED�*�S��m���{c��*�R�}�й�HF�,i)Cc y@��$	�dh�a�Ess�TiEHD}���,=$�U��D("�\�ocթ������0Y̒qW|�NK��Ÿ��9W���*�щ�iD�������������a�GC(s��ڎ��s�s�=!
�4�
������?��$9�CA3s��{o�\k�j4��F�z ȧ!)J�4O�����7�t�̓D-Ԑ7,D�n�Z]]]U�g�%"��l>�{D�\�:�	�4�2���Ŗ���,�Κ���\l�9$G�އ�2.�dN�=�-% (+�����Sb�X�D�Ր�M[0Þ�XA"j9%r+t�)]��T�K��/O��]��d�\2cp�4�[�r~�z׊t��RpT�:�E�G�A�& �T0U @D3-��t*�p[*�󬖢WU@ۿ2���k�Z��(���A��ef�L�;w�����m	 ��&>B������9���޽�o�u�1TU�jr�a��@�/R�1���wV�CZ[n-( ��0<6��Q��I�C�ܳg����??x�0Tn�^���o����O�8+5 ��pBG��<z�H�������m�z5�z���%�֐�uJ�0[b1 TUB�%wf��bF�:*�1Mc�RN�՜Ε����dN�s)���`�/U5���=�G\�m���T۷4��*�~���ֳQU9A,�2�a�e�ttyԶ�یwj�����ԛY����r��(�h�&��@�%	�}��9%f.x�ݸ7��V����U���=�/�n�P##JK�\� d3%Ұ1{��2�B$@Ua��px�Z�ڝM�aC/l�`�,G�`�CTD	]�5>����Qa�UPU/�(�r=��I�q������8�dz����J7�����\,T�P����+EW��e]�y�\�|{��*N�O`���w���Lp��v��Q�%K鑁1ڝ�;����0�m\K����{3ds&�َ��,*�h�F"y�B�L%�2[�އ@ζt�|��"c�J��a�XsFpD�y�D����m��tJ��j�2j�I�B�,��'N�3ZDǨ̆c�P�ґ�s�eX�Z�}ii��g�
Hș�hS�:G��X�f Niݬ��Ƙڶ�m���2�&�V[Ů������1Ʈ�,����.A��*"V�d�w��ca����CL�����f:@�A�Hi?��QKpF|��#�֓������]�cQ�SP$��GܚV�sG���xڬ�� ����jZ�����]�}���q瞯�/�G�UR����>�j�̩�]dAWU�H�9 �&%Iy^��*���P�*��>�./\��GZ�0�u�V��Ӻz�(���@����⼮+O�nVH
�I� �(����-Mi ���[.�uUϪ�y=:Ң���J?��k��t� �������0:.�
f�W��n�� �����?�{�}Ӵ �_�2Yd�
"�r��2��޽���ǜһ�}'T����Wo�j�Z���y��BWN�!���3�2����5E����*�)u�Q�FR.�b �DU]O�:���f��+�P��� 9,�^�n���5h� �����$����g[:>:�=C\OJɨ��mU�:G�����|�Mk [�8��^�s���B��uf0�s�N�$A�H�uvjM}������
�m (�k�`W
���>��Cn�nh�{>f_2/H �z�Z�u�|�kbD/ �_�j�� �F{��a�^!�b$����6���K�9EU��]��"��^���Unx�w�����R� �1���]�9v1v��U��1�̀���
\Js@� ��c.��e���ƃ��C%Ŷ+�d8�f�d�U�L/m�>+���i�"aD�M6�~8h=��j̝P"GV7]������*�#�X�HU�̆�.�2B��p/��{�H0���p0�U6³|@�(1��%���VM<�'�c�Ę���3�z�8�rL���pCoߨ5*�*����ݮ`p8�6ؐ�#S�' pΥ�0��&P�U`R�[���Bq�,E�G��n���ɤF������y׵�Q�11�T̸��8D�7KD$ %(RC-�)�XY={~w2�e[٤6��8]���26%�/�9�%4 ���{��7V�׶��t�"G^���P��Q@e��H�ޣw"�n��\�x畸��y���Ѳ��Ǫ�B[UO��w_�8\�������2UU������kW�N���Î£0�s�g������B"X�^�4����zX�a8�������*
�v]�DuU��l���.w�ܙN�[[[ @H�l���G� �����{��ы/�yk>_7��T�BO}��oz�BSD�j� nD�C�ΆY2���\�|[7A��SP�Q���t]� u=q���Sr7
�� A�4���9z�[o~����ӟ��>l��v1w�uv4���B�!�Y������3�
�[~��R������`Œ蜛Φ��T(���dUѻ�:
x��+�Y%�R��&l�/�H%f�՗U�q`Cs޲dc���a�]!c� ��b�Um� ¹溈QUunH[�Rj�7#�bV�Uj#8�FO���xSQ���^и��ι�BK
��טi�BU]O�I]W`���m����0�H�i��}�"�<��
%�ȜBșT"��(��j
_�!i�5����"�!�"��Γ������ �d�<�=0a�7�s9r��z�_fP��f�5�Ƃi��E������ٿ3��m��w����XJݍ��9�)F���J��H
V^�*ҵ�ڭS��Q��e����p���,��iSh���D���h����d_��7���ϔMv���ǥm2' �j��SJ)�A QWqVD�%�udM1�%
��1vm�Φ�&�p
>�s1v�ρ�z�D�x��T��S�Rg��}�'K���eY'PU��w6=���\�_��l�g&���n�����g��ʡ�TA��ޅ�K"���=4;u��$*�N�
��f���F�!pq~�Z���u��lyo�������Ғ�i�����iڶ=??!t]v���ް��ߛ4 *�(* �
�:d��r&�l�������Po�JD��������L� %�EA5ILM�N�����Y�w�v�U\5���y7G�윐7���{p]G��6̱�¾�V�~�<j��Y?[\>[,�P��w�s
����'��)lm�^7�9�e��#&��K�|�t/O�$������N�y��Q�!�CrHD����:f-��Ȫ�a����ӵ���dG��"��r�z������999�{���奪�t:�洞M���'O�u]7�L������R�x��쒑�^�����Q�x��pE���I(s��f�y��Q�5�������d�i,�zj���L������������x6�����f���������M1r`�2�9��ƎUU@pT	d��sΎ��1;��O&�FO'"BJ�/y1[ǡ#��i���[[[��^��զdv�D9�2�q(R��i��0��f��`PAX��3�����0��%�9�k`��{ʡ��Yp)�xW�r���_��:9�r�~������4 �i>{�:�bJ
cWU��⒈�/��h,��@��z}|xt~vND�������^��4]W�-7nӪd.��W�(
���橷�i���I3c��"[�Ȱ)���	n@cv3k�<�A��FP0RQ���@��7N�X{�h�be�Y1��g��`G�y,{�x�s�(��v�q��ۯ��Ɠ�5D�l=�Ncv�{�28T���|RO+���c�w��Y��u]�Kk�X���I���Z��|{�����Nώ-�>�ڸ!�Xr���*Iae�z2���@څc���Zp�<-;�;�QgK�,%�s ����BJh���rJ2*M��!B5O�b?�9�P ��%9�%Y�ۦqU0���ל �o�$"zבֿ�;7ߚ[��\�y+(x�}p�(`ي�'!\�P:h�;fP�W��/�ؒ=J��ώ�JG�}v���̈�b|뗿���˥�x���u��� �����b�$"0�G}������g�?��p�nJ��2tUe��( �%ؚR�L��9���1{Q`逐�d3ԁ�욒<��@(f% "")��*�rn&o	[���[�=ٿ��7�rg{/��ׂ^! ��&�$� |�(�(Q�`�3�Ζʫĭ�ۮv�[��j�X6h�i�V�Sr�uJ 0Q��G�'eicZ#6Z���WK�����t2UՔ�8�"
�5��-��bLRH��Kf�)'0|l�����ؕONN././//�u�������d2�ϡ�.Ʀi����f�|���b��l��w>����ậ���+�ע����M6����ԓl~�oQT��2�?<�ܳ�ƫ#�G���W���O��pxxجKG6���� ��-�DT�TD�+��T2��u�TU��u���m$tU�ȑ(#����Vډ�Ol)XU�((���{��Yä'�~��&f.3� �F%:�z�d��B�܀a_}s�Ύ�l�wW�{�J��r�|a�0>�Ѯ�EBY��X���@X`3���C릹|�4������KPp���) 0��@�� J亶���o��]�t�h�aJL�Ddv��Ā���[��y��QPoD ֡9���Ҕ��=�c�*"�1n6��\�l�io� *�vբV5�	 bT��L�B+�M@�Mg��NЌA&��^��J�Wd������2^���ҶM�
�m�Y��2�����Qr�'"���|5˨�bO]��{�}��S\.�̜bBX��,|.A����a�|ӴGG��������⬋�h����tIH='��z�=Zh iCr��sp]���N����=$it, (9?\'� ֘�6�����C	�[�akKi�4���j�%X�A	��B��ᆀ*��������e�b�	����s�!�eN ��^�J�sJ�SU׵5Ή1ٟ�y6( HJ�zʸ��x���œ-���;r�l�E�!ш��_*�-�(�����''U]Ǯk۶����]�}J)��DR�I�� PWU]�1���KT��B��frDYR�	��������A�Pq`���r��֜�@��y@�ʒ� �����<{:�dۘP},LU�L�����쓔��{?e����rQ@�9����I��Cl�Ҥ�&�,��ĴnBB�$L.�O��&3���]\��Ô�wϴu�!ъ���[�P´�l�������kۻ���{<�ˀd�b>��#�$
�
�R\�_
�}�;�A.]�c�sR����`�kU��5<;;۞o��Ϊ����r�P P�L'�
�M&�Au$=�շ:( ��U��@A��}}��XS� _z7f���_n�������-�!����Z�v�4~�a��6�o��ma�Z��m�f���L��
0�L���ء�iS��'&y����� ag�����J �nb�j�i4�AV����uL��AJ n#�23vs�;�5"f��9ڰ'E1W6�GI��e:Jz��m&�M�e�4%�����5%z�X�5(���ȧݼ�BJI
�f��v�0W��>a*\��e�Y���i��E�@U�vc�d�a�*�;&n Hd����Z�K�KGQH7���U*�8���B}�$�Z�YD���d�%�Ģ����P�b_��Ðs�n1+����?X�x2�bsL�iA�br�,A�Q��Xr�l��W �g��J���A�W8'��GiX,"Ů}�⹪JUi����?�oo�(8"�>x+vRT�ԟ&��R����6�2���tg�S4kV�l͍`,�� � *�*��,	nx�͓hm�7����c� Y�I��������l�K)� "�*��r:�~Y;��3�b|@V,�r�i�� ^��af2zwFD��>��L��
H���P�Z�L� �䡏�ы��R��eo)[�HВ�pS���i�{�"��R$$������ �y��,g����w�**p�	��VE�R��o�E�<9WU�d���h�|��&h6N�����䪼�6<@�Kq��b^ a>�XgzĤ���]� ���(d�PBQ�1�rp�fOD�����h�X+V���PϪɤ�A;��tF�$檕�z�}@ _9D�jR�s��	xIB,�����_pۨ���݆�㼏�Q��B�<��l�����	*U��Y4�"0���\�ZX=�hW���/z���~�|�ч �'�	(���ά�.� �E��2p��򩪪��(�}��7ȝ�e�?���[�?����< �(1d�l��<������W7�l��D��Y$ճ�3rD��D.[o7�{U%��I��D�)�̛���ϕal,�gaLH [��lf�ڤ���D�w7-�9Rx�L�UU����u�
��}�fVK�r]�!���������53��TU��f
���g Fq�~���R�φ�FܜG8.��tH � 	5wT�ꦔ��KF��A1[,aN�:v`z�fPJ	Y��8�P�;ggMs��C)��y'J]ۚ��V���@{tO�!�W��{YO��˼26o��(��}�7 �O#���l?�t�1g&4�a΢sVAc���瑗��2���@�B.2����ε���Z��rT6�/�g����\���ʼ�#�����>�E�`���,�{/�޻�j��ޓ��ij�D�Q�����!���1&��N��i������Xz`XJ�f�9�uE �F�p�PAS�� ��"[b ��l��CX�ڃ��Z��3}�-8g��ae�`�pj�I�s�k$�3���'�-�2�Č ��}@D�Sӵ��=���9�%ܔ�H�Hc��P� �R!8�� �M�m�B��?EQ*��u�K^i(d�<?�$�0���#Qv��6�0� 7�WKɹ��Jz�`��DT��SJHdmE��E[���5VAD"3Q"r�7C�D����/ �j&���L�Һ�j��"�}㢁K��<�xƹ1�S�lՑq�j�DE	[r���� �:'�j�.����W�S�3��W���	+Ě|��vn����J�R9��y�	z�a�|�T9�^��E�
�!�fs��w�&D������(Y��4�T�t��Y�T�P�8醫�$���ca,c��\׵T� �3�&(Qt�Ox�����Up���_�����͆�#�?��Y{��)�\I$�I��c��%D�ީ\�F/7W#�UNI ڶ���]Dbe���W�O���4ms��]D\�V���� B���\ei/���D�+���պk[��|�:�c��_)��Q�@����]�7�ndf�,s\�0]Yč-9��6hq3���͛!� c�R��z��
�Σ�	��Ḭ��EZH�L�Le�������l�H��QФŜ32f̝w����'U1ũ�8$a+܎t��3� �27BR2>'��,ƍ��>��P!����4QB�¸g&�b���-�ws�s�����s7 �mz 7�{-��+���X�_��-�to� l�:�b��,�r�G,ʨ�H���p�edbndt!����z�&�*T��RL�@A:�Ԩ`�
d55
�}��>�X:���j\=F��)�3%�z�0#�,"�n�"�gr#O;���c��
��ODA��� ��e�*v���`�VJ�RG�*�T�9�%3[][GH�@$u]�"9O���S�g7jXl��CP2��p%�LI�E��k>*"��EN�Z�s�n���[�\���X=���7K	-�tػ� ZBc�$  ����J�b,�T�8�}9�hLQ�?��
6BEÆ(��׎�?����Mi���UWp �g^u����h	<e�j�3�8o#�۞0��U!f�����dr��ĕ��H�W
���`�:E��UD�PO|��j�VЀT��#���(�E�^�����N!*f�$D���:��g��y�)�r+[M��=
48$.H�e:�Ҧ��<  ��8ׅ��N5��� �u�C$6�(�| �.vUU�����C���ȫGc<�́����3W&	������V1��lTQ�v��QX�v��P �\-���1�!�
)%k�b\!1��t:�LD�%UU��juq�888��fu]�mcDD�*�(�[��NɉY��s�dj�g�6�qDUU9�`�wS�a.5��A�񻡍F�'!��9�(ja)"��)Q��](�GD�(Ho3Aݕ���ӣq���G�"�B�=Ȩbx����^,7�qƼ����HRҾ���p*�[J��X��3�M����+�R��l9Hm�C�����ߎg�!�''��$���h��jl ��AR�@ئ�J�E8V��&�mW�_h�3�IWs΋����Z�3�Ϙ*��4������I^����~ ��'��u�H��|SUU��(��`�ح��yQ!�P$1�0vqRUFbeu#�y��D���{?Fu�x+Z�{�Cmz�HBb����G薅Cdfkdi$)��S��+�>(�"d�����4���(�����Mh�7�����(xc��ވ�xf�Ng�9#�N��B!� ��@�z��H ���p��j�$�h�^��5Qu�g�G�T�~!pP�,��q7�j�W�Ĝ��:��<yK �o}�_�e�E0s׶։�7�ԚA�Za�Lܙ�G��[e�px:!�7k�jM�p�0J�I����X�z�'MPZ �
��|�2*���4��+
9J>��> ��f٪��I����b%U�D��!�%��2�xO�
M +秈Aq�pBX#�<MM��N�j������WJދq(�!(sE�E;�]��9�;����ǩ��+^��6l�k[&�,���m��ˣ�yI�s�0d6Z@�N���]�p6��J۵6�vz�r�5� �����.�-�2�����9WՕeɌ�D���(g^�vؐ�����ls�GK�0�+�\�j��Vԍ׆���RT(B 6���"��o~���nӬ/�������_���'OM)9?4�4���,<P[��H�n��t:�N���R���pn�� @䪺�ͦι�mW�ul۪���ZZD�@���=�*��n�W(s���� �����3����Ï�{L��"��j#��??vl�ZB��+��%Ej�f�{��6�1��I��UcJ�JT��ErMA�JBC
�Q����'V����@�f�Z��H��}(�Gk���|����`muF��f�M	1�� fV*���~�������FK�&�E�38����yp����W���y�7n*�̊�
��8���"҇ŝs��y�Q\��λ�EE`�*T)EDg��.�* 5����(�������l�Mɋ�D$��ƞ�Z�:b����	%r��Y����å��)̩0?�Ȓ%6$jέK����{_�u%�,(��m)�7T�%�\ɧ�p���j��۬�j��Ue�!E��ANL�|� _!wQ�]2�g��mP眒��Vm���X�4���@p���{K��N5���u�=q��w�޷��A@J۝�$L��&�h2� @�4`t$f\��.Z�Ͷ�L�8�J�}U���;�tjo�L�� �7{o��P�H-mf�C�%�I2����X�������i�A!�p�@�Б� k*���x!��Pfp�HE�$�
d��ą
�����M�f�\5a��$��bpXM�Sv���8u�m�o�O���9!ze���n���:��K�f��W�����W�����m��Wo�����7�|�
�|pqq1�N����#�p�2��<k��1aa��v�>�ͭd`�ٖ}6�!�e��7zZ+���1B"�H)m��^��
T�,����E̓��	?a�Syӥ���k��x���Ͼ���+����k�9��
�3��P��b?M���󝝝�dbX�y��24Vy7�?�ւu]#�j�Z�V�Q�Yr`G5�_9t�_���x��<�e@�X�"�TX�K������8�	)JR������J�Zg��Fv𰽮�v�/���h@�B�����=�UOZqh�n�*������3㈮u|Â�� z캺��P#��"s�I��Uo��=+�9
p�����<ͳ�gJ�w��j:� AT�!G37,�6�)����Em� �f���" j1H�0\?w4(]�d�S|�_���		PD{�q�ԩjl�8�~�0(���B�Ѻ�^^^R�Ʉc�<:)�MD�X��*�}���Q�ln�>�� XXF�03�s�4kg,_ڜ`�J�q�2���7�(���m!�v�j��e�8����ӊ9ILY_�X��5���1�. |�R�u%Ő�
Lz��,治��+��x�,����"J}ҲX?uBCS;I�V1c�mW�2Y���2��5��̪�D�TA�y_U�*�<*����>Y;$ O�9R��P�r�s�����n���y竪�o�c�qw6���.//g[��tvzzvtt�8�J��K��W�c�O�M�s���I�s[�/� 5��0���vD#�	p�Y�7]j`@�:�Ɂ8u ����q(eͫ��E��23a:u�����D! (*�-%:�@���S����U�A�Tf�M��8�8�P+D�Ȣ�)��R�K���J�Ɍs�p\��8����t��vd���T�����o̦S¿�W�ף�����j�z�o~�;������{���1$��㽷S��)eIg�>�����KC1�������5�o}$TD��
�AR޴=��PV*<� �r )+SnU��MQ�Z�Pv9����G)4&K�F�կ~�������{w�������}�vC)�ᲅlo������je�en����h%e���ܻP��R�6,\��"��V0D!T��H2�qc� S>Ho��r *M�_��NP5�dl����nZ7̆���/2���M˸ᡳ*�l��F����ۙ
�xU���y@�������{��
՝�wꪾ����^<���7�Q���|��'��˫m�]��~#�P��P�4WF�ʬݳ<�Fj�A��c��d����i��~�
��c�h�����xao�`�@�
ˡ�А!mjb�T @��#�75U���6 (X���l�|�м��J���m�3Y��^��㉲O��#$Oa未��~�K�l��u�����i۶)%�I�`=�Â�g����$��E��B� mۘ��k0X���Z�ͯS\H#уbA*���so���s��$�
����h�9�⦔��T[α��v'5C���T1�ʚ�'f��UUE�I'%���X��U1��"��Bp�sde�l���Pt�@�	B1�OQQ� R�h�HX�<KU%%B&	SJ1F5��f�f%��<E�"vf�y%�����{H1޽s�ѣG��ǻ�;������b�8:<tν�������8mDg"Z!�L#R aNCUͶ���u:��m׶�z�x?���C豴���#E�!���>��c7W��@5X��ٝ�̙�GVD�"`Hl�2#�(y�8�Ȥ�� ��@Q�%���[D �5��� ��$A�
�&
I�0�8U��D����\y?�r��\y���۰�tx��b����
��c�ʇU)#����pp���g�=���w�ܙL&|��a�}[-�����ܽ{�����N�...RJ����~�Mf>::Z.WrMqCs�"<C髪M���$�
 ��ɲysCU�Eͫ��$�
�Q��T��3c3��XK7q�B�<����_��_�/��|����������g��rZOl��)��*Bjck0�sn�46�>B��\.���ݻsg�@XV��b�p�Ea� ����)9b��}��뺶i5g�;�\v���=^�b��w@vc�u氎��f������똓�I��/f�w:$W�������S�[��m�����_���[��o�!�U]9r�{�9���=�;�Ɨ���OON��s��^j�aggg6�u]�u����� -./۶uޫ��ۀ[_9j�F�TAW�n��u��f�~��/�����06Nu'c����Lr�ȡ(+�2���r}��i��Z����S��s�F2�ڊ��ߌ���o�M�(W�d{F1��fP�'�7��ͣ�����;w�N'��ˋ�by����?��ӧ_��׿�����O?}�R4�M����������k� ��=��femq��LXa��y|���^Tr�byc��hƥEKR2� ��A����(�!Q!���ڔbN�,9� �7�1o�9�)%��t2�b]O�c�" ��h����k:��ABL���wL>E��؀ 1�d  �9��`|�TZ�Y��x+��*BUTp�@Q-K�@;�瑙�}��x	sQ��k�%$}�J�D$%�a�=�V �0�N����;w�W�����֫�RJ�h;D��&f���H��L����w~�?�`ow���l2�<~���w���o�^.W�<('z�����Z�����7vǾ��n�+U+�̖�u/��5��|�ՠ̆�>�1��>�qT�-�{�J�G���M��
b�l���AP#oA�H���8H���O�Q� �e�K�?�����n�w&�#V�+&����_�z��㏟L�z2���ڦi꺚�fgggX�`�{* �0WU�ַ���u]�������ɓ������ӧO��_�c2��R�A�B>����x����&k\�y�B}������N��ri���\E��I�H<�C���Z��}S��� �)U���Α;=9��_��k���[]�U���nmo����g��j�Z�VUU���w~6�-�}׵ggg���u][�6m]�|�;�Q��c\�V�����ȋd8�S�;�����˙z�%kCGcG�UTXbbP��׾�G��?Z7���}�!#�@TZ�UuN�a�7�m���+S�9�Gd�[	 ���^}s{[�ͦ�ߟoo����د����|N�"Ҷ����6�.�g�P�sp�淾5����ϛ���۳ �s.v���������pAAn���(���
0�9C	 ��ꯍ��������B�8{�bN���Fh[ ���/2	��G�6���x��z;@@��b����C!㑈H
@(��1�I-��y��j�(�������_�׿��~��/_<����׾������r����Ͼ���.���CfQ�Z����Çf��G}|	�w�ޱ^֎���L�-����J1��ei>�!�u���0�WLo/�-�+j-*!���[�e�7��C]W�hR�Z�&���H.��=;b����� �	@].��X���7�"�1�:-%X*�e�=
���'W;Bd�"��U�0"y_,54H�p�g^V�b�؏���`o�TԾ<"�oY�����L��:
�,�{Ǩ_!"*%}���L�qP������R~�9�bPս��G�^S������U�Ng�����>n��{G��)��������S�җ���7�����7M��������]�ϟvrrz}]�p9Eu�7YB����v�M�����䒷�7���66��"c�F�>#Tl��u��V������:�4*�����쟍 I! KW`�@��P�=iO�I�)��a  %ET����@ny�WK��H�*�$6�0��N1?~��ٳg����7ި'�G}���s��ݧ�>],Pϳ=����$N[��޽{��/��_2���G�����r�^Q۶M�d)�ϞX���FBuW^|��6�w�
�#�N x$u����UTv��?~�u��'OC��|��ｻ\^������>}v|r����w�|��O>��ѣG_��W�?������o|�������t2���|����w���ݝN������T���,�\J�gRk6����k������ɓ���H��z�=���sU�b�GGG<�kc�µ7^}66���snk>�N���b�Xpa�+~B�f�f��4;S�%��sB@A �_��?�����O��v�]��|ƹՍ!�Y�o���d)�h�r`�|��3`�X2�f�F@�S��-�-o��!\���k���s�_���|~q�^��ݻ���gg�9r�umJ,̉��s����ϟ�ms��H D5����w���/^❃��?�L�]�`��ŋ���ω�_{�q�l��W`�wچE��	U ����~�n�(��a�5���MfǌUPБU,!Qn���r�Z��Q�������U����.g�Z� 	�� ֒�P��c�-�k踪:��ݻWU��uUM�SB��f��G}t�ν�� ��Я�"N��o�[>��\�|y���|�G?��/���tzyy�^��kZ3檪B���"g59LWߙ��_�T��)P����O3ق"���.���� Z�uUUV#a5�"l)��`<� �,)Ŷm�f�v�RQ�*1�㓣���`ݫ���ڮk;�8�Նb��0<�ID��@�yg�?�h\USL�
�
5s�a9睇̨ F�Z�qʶ���X��P߿j��-�����������Q�i�v��͌�	��>�MD��Dxqqqxx�����×;;;u=i�f6���vηmg�7�To�}�s
*�DT������|����Gm������{�k�h��r ۮ\�w����\��ƻ�^�}S���T��ρ�8���ȠE?��S����["�����MBF4�6S���s(�V��)d���>�����^`��$�a�l*@4�GHΥ���{��d:=??�����'O�|���ۿ����NU�������@����*�ψ�V(vqyѴ".�Kf�{�����?��?���?],ƶ��1�R�0���k&��o�"�
��7���?��?=;;�8?���O�����/�����ɣ��������������O���o���o�������?������G}��7�����������������������'o��{������FNgg'G�ǚ�)���е�ֽ��}�k[[[���1��zm�
M"[-���������^J�X,n��E���r�������>�d&(�S����PN��zU����@�ª�����O��'?�'?��i����i�ݿ������s��{_a(���'h)b5���bV�$<���-�H��⨤��{�Q�$�P���`F	y4�R�)bD
�p�yX.�Ώ�����../�������m��t������u�4GG�m���,O��q�m۶iS���b>�϶����O���z�����2N)B�n��]F�hE�}Y�wH����j������7\���y�J1�zs���G���}�v)��v�M�L�M=#�)1����J,��@���O1n��̨d�dT,���:v�WA#�����˗/�|�͘��w߭�J	���t:��j�\�����5�g�=[����lB��Ǐ�����O����G���7��Ώ�����_��Z����ȹ,
�|�u%��*�]G��.�fjuL@�H�:�,�|8�ou]��1NiY3)%���s��YwB-J.w�Q$�S�)�*Ly"�!x���]S�]���}��@c�r�}JI*��B@P"t�b��F�U����'@����.8Q���X���m��b���Rs ~6��M��l��W�D�dX[��5��-�:K}��
�ڶ��o�~뭷��ϖ��d2��j2��f��#¶mU��j��A"a6��k;,�����?����������)ŗ/_�a����XQ�2,���	P5�@�@�&�#)v�u[_1(�2"׸�b����2g���5��~U+���z�����-�Q�4 ��2W��ڕ%�(]o�iC��ڨ��� "�α�����l{{{�Z�V��tM�loo�um��ж-T�.d�@β[R�����'�|r�޽���'�gg���_���Y����կ�������4xђi���d�����zad�^Rp�""o�	"�J��R������7�������޾���>x���CPI)޹{���#$���?�ߣ潝�G�;�������!�w��Ǐ�%�p�\��J��e6��f����_����٧�0�|0����v�w���j�
!���i7�f�R��s��U]���ηfm9F2��?u<υPs��`��^��  @�����?�����x:���KD�M��G̜��_��Ó�hğ�.��&��O�}5Z��,��4'tE������� �������?�� 2�4g����CB�f�~��S��u�������b�T��lvpp�5��x��fUb5��}p.�i��H�w<[o�c�*�fQ�V��6����A�M�M�����Į=R��=j�W��{����|�ϙ�}]�7�9��󇝝�;�DU�'��z|���������b�:��D�V��ښ�b�Z�L�R�����f'����O�:@<1�ڼ�|=�j�����ЬM��"�0��[27�!�8�B��;0�<d�]c�u�Q���h�I��'�YFt�L!�A n¶���������1^��^ռC4����C$b~��jeշ1po�SLB"�R������8:������RP#�=�d-�� t��=q�.�"�o)%���;6������S�� Lc�1_�_=-���� uI�U����6�S��ݥ�0�eP�GD���g�\N%}� ���W��1�������p�a��KG�h��Q�SeEmMٲ���6Xլ�^�I�n�FK��)�+�q�+����F?�N��$ *#��J�s҈��|��^�A-}�ݦ�LwT}�Mj�����l�(�8� ��,2#w\[���t^��2�3�NC^Ad_`�\�`�I�m�dA/h�Au\1���A����ZdѮ5����,׊_1s����>�(e-��2W��~l=}�2\���%M�!�,�¨���-k�4��w?d1p�_�9�xf�c����9WΧҳ:Z�q��t�w�f�5����7SP캶3&�d�����Ƀq���|��x�^Ϊ�g��yaF����vkSS[�y�E�o�}��^ͬ�,�:�a?���Gm����.G@�Z w.Q(r4P��'ş��5X>����0 R#|P�Y�۸����ۻUOeo`u"��sɷ��dB:YI�������t��h̪6f"��S?�������*���1he~w���+��0פ&���l�|�m0<u�T����On$�Y���ª/��,�s�+΄����E!��F�=pg�d�̚w����lT4�VN:��M#m���:�a�%W�����j��u�G:m�S_��1F��]]�?��?��	���#�
	'���b�x�W���A^�������Zͭ�t5�v�\N��Bߍq�*�8��橽FП-+��Jr��d�f
�%�E'$t9��v��S��/\�/366����(��~e��3O%�D^'�cd��������}�����/�Q����/Њ�>R>'v�ݟ�q �>�Y�s1��r,ab˝ʌ�;�J*�����Qw{b���+&u=>�n�t�Q���_J�~�ʽ n�TE�{<9@3oN5Ƅ&/oM�3K�t�o'Q�ǜ~�oC}��	[�~;9̐�ſ�}s5q���t3#Jt�E@g9w&��W�5C_����l����/B!�K,sj���ّ*�f�f=>��|�O���4�q������v��7�N�H�6t6/'G������p���q��mp(��y������Nň���a�՜���4�B��gN���W��lLIdQ�sIL�~fpaz|���Ll�v����5��u��|�����������5�Y���&�P@<�.�M/Z�<QD�j��kkla4 �ID}����C7L#SZ� �e�W���	��_��&mCl��\�f�|���bD���;��;q����7����{�+cp�,��mm�]1�����}�����R������Y������ν;;;��;8������Ǔ��E��������as޾a܀N�I��Go�ޣ/��5���iH�c�L������PӢ���wJ^�M|q~�q?���� ͋ؒ ���M����IP�1��|�	���c��f���* ��B���7�/�gS����r�'�向^�2[}��дB.,��}SI��ZE�/��J$��ڻ1\�%	�*^�}��_�:ӿxA6�omFǙ!���ǫ��zA����bk��R̹�u��:�/��4 �|9�(�I��qb
a���I��>E��7Yy��$�HKI�":�����fL���Cp��k�����|�6U������x0�����]=���.�֨�((���l��=��Gљ,������D�V�)A�d��(&---!с��z����\���ViIcs�{Ѧk�A�����ͭ��C�Nlx4osab۰6a�V��
�o�H��ٍ-p��#{�Kt�ݺB��<�c���1è�!�J���_۵�Er�C�̃��&��z�w$|���o��0���r?���Cv�I�mΨ�#z�T��W�'%5K���Q�;C�ܾF���Xm---F�P#����6A!��=۬>�`�jSs�����鵃=7t�N�4�^�y=���4�W�6𪫫K_o$×r�����!�]]]�����j�-�k�s �j6����P�����$�~驰y����O��|�Fam�@>r{g��)(N����؅U7���G��b�|J.�HI3�F! ��h���F��UZNb��P��7���J�����ڽ���Ԫ�V�)��B���.p�����t��k;)��att61��v�.�-�0�J�MNN�''�� �zf�0�3Tn$O���+u�I%%%�`Yn�:Q��'�`�j�Н�^o=&�w�YvfS#d��P����n�ӥ<��/���~:�m,���-H���D0*�ǘ��Z����{wAc���[T�< ��E�7)�Z\e��O�)����wYξ)9�鸜�Pe���f��tx��B��_ ���1ra�#��^ha�]�w�V����d����@�4e+V���EwB}�,����eI\@�� �8��k��СI���L��k�z��Z!�1��~�~�2y\�Y���ov��P`@�������kدa�� sg�V�������]���;*i��b���xx���^?����;}n�Hp{ɰp���w�b�8�KGé��Jh��پ�S�k��\hQ�C]W��RR?���-��|���T���+ӓ}c+t0;��|(m�v��j����z8z>��~���"������4���VX�-�G��q�X���l�=�{�@��B�z�6׍��#H����M���H��Z8< ���ډ�Bם��]"�D>?3��d@x���ot�__[3Ӛ�>:�)�������X�������W�آ_���f���eA�9������J���vQe)��S���~/��7#��j����b��̾]#<E�M�� �&{c�����;��Cv5�w){�ǭRG�X..��-c"��zE��lÈCP�q{�{D�g���6�� ��21&��v?>��R�lX!l0��oi�	����̰h�q��HV&F��;���3���w�~�'/���".�mi����~<�$����o�GN�h�.����5x��\5���x�g��sS�r�!����j�'I�+�B='�순���U���r`�\�����_R=Zx�.%�%�-�\��DX�l�V s����6�'y����U�_
�O����efE�uؿ���5e}�r��ʣ#���ҁ�����^��v�J��P*sΥv/����ɉ��^�x8�;8��S�Jߠ�*U��0!�̒.˶~T�\�E�ORL����*�R�N�sE��^h��x�^��JHh��#VDP�-o��#Qh�0r��-Jq��0�eQ.���e��yoZ�l����Y��UG�<(kl{�]kw�����J�P����w���<]k34�@ज़©�(�2�@ ��Ƽ../3���ow{{7O��o��:Os���{��:/���pv����Ԭ'�H^�l�I��b�!/������q��[D���4�Y����~8ͫ??^�R� c�8�`&Je+�=i�!�����+��Yb�aOl�������j��b�Z��u{�]!��nFL]+��T�׮���¥ir���N�Qe��)2n<euA��c��˘�\�����"���.��O'؃2�y"<���Y�ſӤ5�d1��,��� {mH�<M]�~*-6�Jg�GP�S� hC���Mx����}}��G�˞�z�v�`_��8b���F��lR���n�q�|��l6�^���'c:��'&&�ȷP?�
�*�tX[��t���k���,>ӷ0Ee�F)���^��BF��kɐ��������s=q���S���	�����s�;�w��}�K�I+m<�Ku����C�تh��
�"��df�{�v�F��O���H&�GYF^�ю��*�w���gYi��/�sV�F�W��7H��^�d�`��%�D��(����j(�/����o����Zx|�/x:���5�:yzz.w>�Տ!��CCC������� v��F����Sv@p�}~%�/F_����.��K�(��<���֌��R��Dq�3�@�"���㥍^ۛ@пDG2K��%?/�i,�b��y��#r	�48ۢ���������؝����V�k񯃶Ɯ��bťUodaxzӋ9��VM*�}���ܠ8�p�D��d�.)�+��(����58�*j(&9,"˨�.:!����7��Wߥ�V������Ey��\�S�9#M��Q�7͏�whV�%U��f]���ObM�Ip��V#s��_ҹ4�k���Z�m��æ-����!2���u�J����֫�d�ߚ�L{���"��VÔ�_��l|�BN���.���[�����k9�j�e�hmf��p���U�Ŕ`[	"��T�<<m�O�C�"m��ⴢ�YX�Ծo�	��D�ݙ�@;[�m4e:	�>�>�������~�.Z���X�ß�F=������`��2Y���c�NחI��m���x�K�>�1��������7�V*�q�Z����������W����n�31{*9�^<����A��&����K����;�Jx!���z���瀣�ۘ^3{{6؈����o4Ԣ�����p!-<`�RW�Q���V�NyH-aY��qMR�Mn�Ko���i`�/>r�&��Q_�ۑ*�-���b�I�=7U[m��`/6p������Z������lTܐŷ3������5�tr�YQL�`گ����eA,����H��1��i�Z�p���l��DƟ�V��i��h�b��*\��w�NO���s�R������9���)sz@M#���m���K�n߫����U�|�grs���{{���u��{��pf�t�ߘSZ��o�����--RR��󇇇�ѩ��?�V�t��zmӬn��ޔj{sg��l���Z��X;y~����J�:gy�DO�1nZ��=��ࢴ���B5=2?w,�>W}���C�@�4q��;֒F��oXJ��?�ϗ�OOi���EC�Y��\����Fh���e#�l�_�i@�qm4M������Һ���^�����Ϋ^ދC�EіPО^/�=�֖�f� -��]���Ã&���d�x��ôs�-�\��1<^���<}�������%��׫�h���������`�>[��l�,K��d����P�l��7u)����ltv0�JC��0��^] :EEEqz�''�;n��y1jH���z��?9+�=I����5�3��4��X�:Q�m�w��kN��>oXO����^�:��&���vG��H�~�{�j��h�=���0)�ɦܔY<��s=E�(�qY,t#�۳�fE��x�7��1A��Y[��q;N_�k��B$?������=X�~:�
:ޟ���3u�þ_��,�׈�r�j*h<�9YߥM�7���V�р��[1C�?�۩�w݇��1dg�52Cı�����S���sk1�Ϻ�/���j��v�6���^0仠�����NO�{=���%{�s ��:�c��iM͵�ؒm�ۼo�N~T���Ĵ�P9&Fz�x�S�ɻߜ.���<��W)
��F����gc�[��Dd�?qM�G�0>�AWt����4k�GbN;�^_��^;��ʩLײ[`��'���v�?cjt��]?9I�eEIp��S���R�>��m�ٷ���YN�̤q5C_(����|�\��.����:��l"�!��	orDÈ�����naq���U�h���$�m�V}����3��f��j�k���iv�H#�_]�j��a�3~B�=єP�$���6�wR�y>~ǱK�btA�
��
��V�ـS�Q[�1�J�����7�U2�M�uo3�%3\�r�ʊw��m5�b}��{/��N�3��MHZ�e�K���k.a�����C�c�g��� 
M��M�l+�k�5��v��y��)sW(��r���>����-돎677Khֶ��g��2K{��""x��;E�ws�[Z��<n=z��Ld;
���G\||�%���'��7���y�&8\0�Q���T����{{���dNN��y��G\�й]������
a2��WS[|̀�0�(m���%8�7�4�(�NƆ0j�E[�'	�<��^=�]}Z(������B��sj_�_CVA8C�fOtK�;+w�`�J�͆�f~0�Q7͎�h=�΂6E���sI�-�T����y;׻� \�
%/Ƭ��p�I�҇��K>V6s%'�$�Z[[K-�"�U�KL��~�(������xu5��^�x���L�q'�8��f,��:��B�����XV2<��T��ʎ �,:q���<V��� ��Tm_,y=��$������G���1��^���y����n��o�ֻ���RXj��l���7I��N�3|�]BJS��v�W�:��߃o�Dg/�@�iO��=�L��-�"�j^��;�au��
3-`�@2���l�v���$�'/��ƕ����#W�E�C���#�ښ�o��t��t���wt��Ŵ�$jC8HCȘ���$�YT�����}Z�)r�DyB��ٶd� �$�򽮳�Ƣ�xRJ#��XLJIW�"`�&��<s����_��6���d/m��^(�b�]�SDZzh�a�Һ��i@�� �Ez�<�G/	�Viݏ&�0����������>G��Wp�=�Ӎ�d������e&����j�s[n�?�vu��A��C�xt=(��N���a��ꀇ����KO//D��^����X�!a��+Ye?��_���.��p�׈��}�c��N�h�ړ��Em�Yc����8N-W�Iǯ�}[O�B��⚔}w��^�la�7�����:sޕvW:�4`�������&�_e"�rj*ڪ�-�r���09@B����������?u�g� ��>Be^���.�g012���y�D@"��l�+g��o�"O���"#�t��,?I�bRK�d�Y䭱��h�j�=��!����:�e]�Ǳ�~7k%ԫzo.ζ�F��J^X�����W#m2?Ԓ�}��`ƾ�5J9�O�Ґ�B���G�_pZ�#�%���Rok/�|2ji���W�kL��!�f��˹��y���v�������|��;$.��r��F_�{���;3J�U��@��V��j�k����q�SXUUռ.��j{��vD<��>'{!�[U���w,�!�zL��ٽ�׫U:��~�MU��VnVL����A�+Hx���|��?Z���|Q��4�<�1o^ ��:�7hj*G�W �����!uZ#)��i�w4�o3��s֦�m)�ɿ��xCE��2]H��",;����	8	l>x|��E�� �l���	=��+��\�O�d	��Jg�t��" e��ou&��]�xJ���۫c�_CO�H����I�[<�+H���I$m�$�p���f��4��D���~z��{�����O�L��4�.��]J��O�`Z�뢭?k#E�k��_����iȉ��y�%v@$rr��an/�i���O*`����mq���\J�_Q�-R��m�o�Q��[O�;w�*��t���9�|��M�X�%Ƶ܏ ����^����)"�ۋ`QDA	��3D���V�0��^,��+�~S�ߖ��uƔ�������f6�\���}ii��2u�Pj��Ґc�Ϊ��^�ʓH��qP-��=>�S�4��|#��%����Ke��m5K��+ W�R-\�������/��^5&�(&?s�I�6>�M,3�W��0 ��K��e�%`�g	 K2��B�tu5Ȭ��^[�[L\�\m{�:r���� ����F)	�Ed�:�z��������X��>��|ݯR���e\
����xh��wvvG�����'f���ǐ!;ҙ�gV�`,�f��ΊҺz������r*gj��y��Ќ�����ʕ�I�� E���U
+˙��R�N��
fy=�W�Τ�i�P�s�%�fE�I�����73� ��~�����8+�\f�b�&�d���@�!�sr<��b��%�v��P���]Pa���������pt�xi�t�	р�u�U*w4��X���*�� 4
�_'�������	$ؾo))���p���Jw�Ķb�S���+Ӟ�v�`>"Q���-YxQo��m��|K.�Q���+V=��RN4c���W�	�v�;<F(�Mrq>7�L%13ۓ�������Ƚ+�T�MA�:z���ֽ@��������?p!�@t겳ӯ�hƞ�9���8?ˋ�Ẽ��Y+��j0x�5��k���Fz����<==o"�u*6]��xV(��q��T ��/���pIiQ��ǃN��Ry���P�y��D3Uf�Rݜ�����6�t��=f/ߕ�����n���@ ���	{d������M�[Y���!�&@�k���ڗDS��z
/ϩ��U�Y/U�P�q+�����%=�n�v\|=��ktt�dζ��k��ћ�,s�m��Y����,����N���D
�]܂���=�a�cP�Vd��ɐ�2?�����,18�du{��K���'9��#a��B�-:f��z@ ����-^DD��D�BMnN��q�
J�+x_*�O�_�؛�{�fsʥhR�֯�+d'�y�X��%��w�5paD�\�����yn����	ր�^�crqǎB�e��Ix�DJR���nA/���wO\�^��|�f���3ݪR�d���t�٘¦]�UmԐT_'ll"d�)h�f���n���Y��t�"����Mz����ܞ���Wp<�����W���2�6��x�+���#��L�)̬/�܈�����F�g>pmr��&�e"�6��FIw�ߒ&�8�4l����X�����W��GJ����qx��[�) ���C�("�}Ӂ���>�!�g�!�{��[�H�(˸^�[�`䒟�F�����|}�-X��^2��(�=z�<��_LD�����kå u��xFy���ο	�i>��3`�A����w�_�޶�J�E��%צ�Ls�o��L��Z���΁�l^w��$�Ol����;�1���<�>��y���g�Gb]	Lh�X�3^b�$޼4X�D��[�'a������J5! �7#׽�v�Y*l�����]���sv�n����DK(�іrQw���O��+��@q��$���˛6w����af\F����h�toԾ���$֓	uc��1E�����Q������~�?m�_e�Vu(D�(>�x; z	�`T5Sq�Ù��� ��L��}��Q=3TjaG�ڤ��2�9S�=�0��h#'�"m]a�>.g�ਇ����.tV�y��&�l}�H
_��j��� uG���V9,�T~pz-f7�#̈́1�8��g^([���v�Z��;�Jbh��tx'�����s����.Q��7g����M�Y���t�m}���ס���<^��*Y]*s�J\\J�������A������*
�r����-�� L��׵�H�dڲZ������9��5~���B��%%��(>��mG2ns�$�9=�rP!{�v��dc���A�(�faOl����yȪ��@��́o�|��;�[�\'F�)rk9�C� ؽU�͍K�^c�i��f^�5u�-�D�%n�'���gL����\�����޾Ѡz֞��w�|CwXC�TX���Dת�fC��:�S�r��y����}ؕG�ǡ�4�Po*]4��zU��*�0;l�:�X���i�E�����g� 1�+i<MLWL�>�nŵ�T�Z��)�����3p��@������ў��>Q�0SVhx��s�����s�k,O�3��/���f+ L��V��8,�����1r����_o8��}]Sz�#u� �y��o��rZ��������F�P��m��k�����v�o,!��z����N�Is����_�ì
��߂��&��U�y�z�$���!6(4���q�T@f=/�鯁/��e6����y�]����ࠞw�{�n\���ʁ7=�����J\-+��ϣ�Vgq�R�~%���4(�nxdMd�,{*XV�v���h�U�*�$S�XBRxu��>-I-��/܅m�/��	�S�U�/̐f2~�Z�+ᮼ�0"����t���ᔅ������G�AE���~��3��Q��M�DV�ȏ[�ˁ��W�Ǿp��[�����T�	�r�z���E�84P����%�3��}���k�c��Y����J�|���ˤ���HKj#hw���u�h^�f�g0��+���Pn#�?BF�$��8�lZN�E��Y��2�s�ј-��Ȥ2}�륣�򀁢�K�y`8I��N�}��*A� 1Ϗ��x=.��qmF�`��D�5)�*j��yKۭ	gZ���z���x&֞�p�ˏ���|c��^���_Y1m5jp�V�������P �2�����kK���EK����Xphb�d:�����1�,��+迻srssg<������a;�Zj��(
M>������uO�ܦ���~w���2����"��q o���I���w� @H�q�$K��^�	I[h^��$e�R)�Mmx,�\Jr�����S��I,ۓ�j�;�Ok ʾ7��F-���+�J��.��!�w')@Q�-ݽs<����I���J�vjD�#			SI��Yx}y�Ӭoi\NH^n.Sac1 ���p�f��&��`������n����]��`H�%�ﶥo�:jr�D�F[�gҼ�ֺ��0�P�P�c4w5�G��rf�"7����	K�"�*�Hg��)����=5�g}��*ٗ�,�ו?W���.�����ї�L�ُ��0��sߥ&�ąy �/�����]�ě�h�h���/<���v᱘%ȼ���A�4�J9�q	�4��	�.1Wb;�U�a*��.��p6`j�K�nM�y�| ��P�O0u��#�,aNXP�{����& d
�0+�kr�;1iQpȫ3$�Lm��d�ߦW��P+�!�T:򩂠������ ??����Pz:����Wa�����Z�ݴ�-9�;�����Ո�����@X�v��	�q^�5�9��24�i����Q�JQ1gW]�L�cI���>v����:��vZܹ�S�P�1�Fq5X��^׭%"g4����	��ɗ��Wʐ׷���|���l�2*�����Ŷe!�,GG�6��.�,���D](��􏎎�J,>Y?1Up��{rs�^/bf�ГV��-?\4���c��:?�.�3(���맸I�N!!�:���-c�N4�%'��^�v�h3�V�.�Ɖ�ʶ:���i"��{~�Za������,`�.d���=2�IA�+�_�*��J9��3:���Q^̐��v%�Q2u����7T�\2}K��?�v-�!ք���Hp~N�7�~v`ffIE'����>��U���V��1�V[f�N�?��p�en�We:��-��&e�p���c
�ǭ�"�?�o���dN�}��co���9�P�U���X�L�F ��#���ߠ���]4����B������n�����媆o^]��E�Z^�ѽd��ݡס�������<�Hü�>��z��Z����ݱ��5��� EU��kQ�~��oӆ
a���'�����eT���/�/����	t�bs���O/F1�����n���B� �V-)(}�/�>�?b���}6Lit�~0t�P:���� Z�Y�g{������!Jy�\W'fN��u&�e�뙼�w���h�b�������<��n��WEH��|#\�a�[���;ɨ���VQ���<Ux=ӆ%p�EA�`m�5���%]	�Ʌ�eqv�O��p��}�g��	TfS�q�q�.݀�v1�M����d�J�ښ�BYXP����W7�3�R��u���_�6{f^�g��A������2��b6q"�y]�Ds�E�ޔ�	�G6#�a��n���.��=�E����x�1��~g��ǭ���}$�_(�Q))���6'~/�C4�tW����hG�5��<��y��RN_�������8��I�*�|�,��111&�7���i�h�Η�I18��{��K��O!��J���͉���
[��sy�V���)��ZV�Z��|UaiN����ι>+j�s BB
�V~�(p��<������D�W��v� �`Q����6)��}M��[x�   ��+^�1��p���g�K�l��㩆�C�T�_��@z��s~�ې;�����Z�BJJK�s���WQ�A����;���F��V~R� �w��Y�+��3rߵ�������bs׾�:%��K�E"&ٶ�p��@hJ�:�;�8$�g�WJ}���RۃٺS|�0T�������E�@�s�W� h��Ba2�cV���R䴻�E�����o���Ǉ'zi�U�<�����s�,#+�I �O@��~��?�-�a՚�o~�EB$�>_��gS3eW�2�� �=��y�X���(cz��3�e)�^{�vp��^z:զ�Q?�yW�,�l]�r/̥�[�_���� m�(�Gk���#y�3�����E\���w���ln�؜�h�Y�/�G]{]!`���*���1�K[݆�^-�����]	О�Q\��tP�l�~�?+�!$���]�a h.T��F�vV{W�����"|�ފ.QfeFƺ7�V'FJ�
��vf�\155G�����\��v::��7���������y�ҩ<Ca%����E�:�ո�)�����$R�8�ɧbh�,a\j���XI B�ж��
bO�.]m�6�F�7�"jMY֜l�OS<�PD��h+� o�&Nx����㌍ZXt#��qL�=�-�&f��$�����ƕ��4Zz�ʕb'�z8�Qn3�/H"�[2�tN^R�z2y��hڛr�5�?�i�S�qS�<��w�E��N�l%ߏ�z�_>9/�_GBgY���+��`0�GĹ��b&�����Ӌ��|�zRs�W�}�3��,n���0�֫��L݊i�%=��'�.��m4'F�?�<��S&]�Gg�ˀ�J��Ҁ���t�&��/�Tf�&�*j�6lh�lў�j?V���=�[W�j��C�=xE�D���!�HM�,��P*�A"�2�W0�.�R���=x����u9�������6�?���U��K�7�q��������%�¨<�I��W��l���B�#D�5Ʃ�����\����"��Qf�\��L׵TeD?���:jos��|2t��9k��8uٴ:��n�� "�r� *q�t�v�q-�ʢ鬓�����gL>�ne�H+�5^k�:��"��e���E'��jD�a�~���C�k�dZ���i��+�,���)p�~��x�j�$;T�Z�w��\ 䨟Ԡj��Ss-%�ٺ3"01��1�`Y���1�:d�msB#m�t������CVڛ��Ӳ���k �K\�hB�n ��tvyO�!�L���Q�����?dg��)�IZ$usc�����6�/#ۢ��#�]0WM��%Q-R�e�(�Fh�Q�vlC��כ.��ϡ$���e���q-G=���зN#�]Tf����t
�@ �H?�g),��0L��E���+�;���5����
z�"�,,o1���˧-&	ٿ��vW�v����~Ҩ�E_�iH*Y�����T������[4�H�=�⵷���M�����=��k�����b��=E�xj1���������'R6g35��{w[D�A���ʺf��4����3g1�/��qPl�u���nN~�,�OO���:��٢�zs����]8<}�vָ���d�P��5Ś+}v3l��K�?�ȵN� \�,�Ƹ�'��Ou���Kt��k��$'���؜��?�gl�s*�Jj�Q;{����G��h����yc�)�?S�0.����^��1��f�&�_,�0�r ���z}@Y[��r=F�V�|b�m5�yf��[��-`�>��@�;�!�]ӉA��ش��=� �<0������j�޷���K|m�9�����g4��[#~��������5��H&��ݯ>��p�R�?Ǥm���\�D)�3[GI^�5�jŖ������H!�L��y�z���Ď�?���{tL� ڜ(N+:.gs�V�VӜ�)}"g���v��ϵ�f��] '��z�+������<��\���Zks�𧑃=�J�_���)=xaZ"^ک�!Ì�Jfo��H���8�uÁ�9Oǆ�T_Y}ɏ�������ɂx���yz��Gw潁N�.��?͔<ja�[�U�>�}J���e 7��)�W<�!�<:R~kZ��S�m��8��g,I���$�6wC����������V��8���Q�}���;dz�ז�0�\��U3����e��=��MH�K�����Q�?��%\��� %[돇,�5�v-%ބ��*9��&O�M9}j�̀@J&�V�?X��V�L�Tq�H#��h/:#9�~���}FJ_DS��֑��zMY|�e2Rxzu>���P:�}�*�������PQy�8?afei��tk5/jM� �I��;ƥ�3&2��\8,RI c�s�8O�g���4�ʒc#Wl�j7������a\-�	PLZ�b�6D�w>�w2o˜����.?><�=.�3�Q5Wq��o;��Z���Оn����^�O�𝳄��jP��[��,G�m��A��2�d��_�W��Z�߼QѮ��ȍ�M걿}+r��^�n�zdA��*�${ap�@̘y77:�_ٴ��>�f��&Z|�s�\���YZ|;'-GZi��H��¢�=�����A���"�U�������?N�#�+�}CX0̵�\T�O����츔����`�,��o�1��:_ǽ��!�j^2S1�dO����@���֡I���]��ZN�
��$7UL�B(���涮ڈE�՝	�uP���/�Y��W��p*)v���V9��ZqI@ꁵ���?e�)��΢�p�,A�J�w7�d>'��������l�?�@�d��"`�i ���;��'Z�2�_ᇇ��%7�C����ې�;�����HY�vq���6,�;�v��Q���ܻ��2Sױl��<c�zғꇋ��b������<m�/�<}��U�<��T^^����@����z�����n��޳��'�ѦUQ��	R'� ��<��#��3�2P��Ϫ��(�?��j{�7%���[��$����=�)���o��$�L��tO���?�/��ܢ5!t4�����K�b�;.���ڔr[ݱ	�N(*9����0�y��� ��~�:�E.�yd� !��$*5��S������u�����1k�+��Ǟ�H"Y�)�	 >�������ݾ�ʹl2��6�73�f������5E�ki�Fi�m>���PhTQw�k���{Y��:�iP �p�fl�x�Q0-�~��I�6���T����Z>s�`����3󟶦��6G�	��;WR�y8�C��.�ϵ�qP�"u�dO�ǵ���)�بd7s�,5�}��R]�~q��٧A�l(4�is�;�,�Э��cX|��������૽I��F�z���Ԇ��)۫�ۜ�f���*Rs��;���IH�c��ɺfR����1	��|1-�����!�q;3l���/�u�2|T� ��R]4]�B�E�/�zP��d��E�:4ԴW?��Rc744,�6tj�ƪ�p3�3�"cUR.@����i¡�+�nҤw8o1�� ���rr�U���'�K�,4ä#N���������"Ds���Z�������e�T�TX$?��|^����s���U8;�s�n�hk[�,=y�2�7JZ�V4��VB4O3��uyS��3�ῡǘ�[ҏm�E�G&���3{}ϻ�3LPݱA|��*W��^Qa"�� 3���<X�Xܢ����'ul-�����!�i�+q�hs+�ZQ�o;�0G��OW�Δ��?�E�U_�)d�}��4�z���nY�>����g P}��3SQj;� Fٱ�DF���g�A �C�F5�ܟ
��>��
)����oΞ�$�H>�/�5���sd�
�����&�����$��W�M4#	 {1���i��ٳ��6?�l-P�� h@��]�
�8$@aQu>UX����3'f�����q�8Q"E��}U�\�zcK{�=�fs��&
u�U��kˁUP+�$E+�!xOb%D䝧��ds'a���s���*(Q	i�� �yc��q���JbD��>�v�%�&Jʩ�S�)�ضM�+�����V��[(����&�d:�z�
�j���-t^��`�Z�����K�"�#Gf��R��,V��VoA""������W,������_����%���p51?�l��va&S�U(���� �����.�T~��e����Ǫ h7X�J{`�; �s��1����� �yp	]b�j��� ͛��U���R� �~AnL�B��1ۯ�^���7�x&�H�|s��ɨ�Q�{�޽�}���=��ٳ?�h{�}rt�ӿ��w���?����1��i����E4E&Q��g�֔�X{�^eI�`9� "1qp��j :rm�.�rc�xW���u]v?�3G�|ldu9�,g����j:�
�l�5�'��k�n���&��*��O>�\ńfS��y!�7R��.�i����'#j"$H)5�&ƈD�;��Dn�]J͙���u���l��],B�<f�r��1  �����W\��� ƴZ�� ��$I�ȑg��52|ˇ>4m۶�sd!h�6$U��쟪"!s��)-ӛ��l�>& 7��/D$t�ʜɏ`P�o�F:n���є�~�G�N��-(�����y��ۿe��J����7�����8�� ��ҡ����Ech��"b*�K ���q__�|�1����jQדz2!�9(1՜�O �ç
 tm׶���ч}�K�Sս���iV�U�mڏ�||tt����n�v�T��U���^Yq�J�nTf&�yB���0�$Ƚ�9K$@Мu�J�6�@�Re�k������Z<1�0GjۮmCU��jMd AA���5>s1�	�l�ܤRT�
�� Iԁ��keV@r������f�<�.�h1ۼq��D�X�>�`����U�H���X"�s.sVAޯ&���/����.(�e���
�(sJ)5M�����m5�Y�v99	�qd+e0�d�Z��m:"Kɾ�`�� �*���b�]0�1��Yk��~���!D4Im@m"24~lzj��4B�񲙑�K��e,e�$��-.�Z��-�K2���N����i�ߍ&'Z�߃��V���6e4˪�f�(X� zȹ�t6��Ydݶ��(#�^֋��*���u?Q6|*^V��v]��N��?6FJ��Z|�ܐ�ʡ+�oH�P�[������7~��ܹstt��lo/�_��Kl�.q���'���DF�N�l���58��={J5C�uf?���M�Z�:�FO����b�.yc�沍~�L�"�����bl�vw�f�X���턹�;Q1)��������x>{l8'�dy��o�,3`�P�S��8G�j�"
@!G����9��I��<���="3�v�[j�8��P��}������Ό��H���sN���-3#���> 0�Ȫj�
J���"#��̀�0��G��#=��{ ����"3����Df8������4 ��������.]D���gw/_���r��i>�^�?��B'h����.��|9�N�����s)��/G�x��2	���\�a�vk�O,~�5ه?K� x���2f3轫q|*ySG~^�������7.��
{���Dc"I6���}�*>*�48�$Ƭ����XP��� W�����ރ\Cg�`<���7֭w��ϟ��Ld�}m�lG��)�jw��mmH�����~��"$Q9��Wf������bf�˹�rs���Cd"�1�?&�QE��S��0�j 1C�t��ND�I1��=l[W��6\a�D�Q��I�Xqخ�/�ւEDV�b�I�"*�WOB���8�C4���:��d�j1@�����K6�d��b����ifN<���&�	�ע
�BH�f
�L*�\�
��GO��/DU`�?H	v�y\��z{�<�^��>F��P?�:�	JY;�r�<�S���U�}1�˟|����ϋ�&R�)��C�-/����7���������	`�6d6���y ��^z<l�me	�w�P���pcOL�Z�нG!�A!��!�Fo�V�+1�L���ǔ����y�oo=kf{\�2 �r�\O'ǔ�������e�_06s%��b9��tX D�=�h�TT@3�F73&z\N/���ͯ�����~��WD��O?}���_~�%����wU���/O��'3��\�xs �e]�˂��77jv�p�����x겶����z]���XJ���y���㺮����c ! ��k���K�d�>'q9b���.��(�C3xxx|�j=��j��۲Fi�ד����b ��_��'����z`�Y�*�����R\����|zP�ŌsYB�=�,]���Zvi�+���sr�#@��M�$�
�����������!���<<>��߿{www8�^0�3��r��Rt��=?�O�� }b]'����Ld��Gt�h������%0F`Fs�H3�}E\�ht{���3���b�TѾ����@�f{g&�#��#{�n��Yx����"�'��K��'��4�8ð]C�D�k�R�emk�)f*����]K�nbBK"r�,��(*뺨"2Divtj���QL.�33Q!����;���Yj������/g=��=Q h����^� �-s��)K{�\��]��YDD!��~"Lm��tf6�Rx��ޚ�f N� �����p�u�SP.\�s;/˺����+E�1s"��Ä�h�C30ԪH�3�a~"�<�z'(F��vB��\x��]��S������C�qL^�^�va�݌���8c����%S�ˈ�,� f&�"�^|�,*�Z�um��d*�5��4&of.���`,�)�R64���}�'���<�]ӡ>rM&��nf��c�q���."��K��D��n��V��?~�ZN��^�ros7�w}�n�\k�A�6G�{]����"���nno/��{������<�.  	����p�&�w�~@�~��i�)��"� ���o
��Vm�6�n�ŐFܽw�+*J�o߽�ҏ��˗/_�~������7�JS}��1�uY���<��Jol�[�E�>'ȍ�� �s'\���]z*c��hԍ_�H� <'�21j��u�>�f� ����tz��1_��'"G���!t�BXK8�� ����I��
� �F-~�Q�GNLe�\'3a 4P�Z�FP��>���l��S����y�[,g�7�hm�r� ��v�l%��*uފ>~�km��\x>̷���z����-S��$T��#����oޘ��xT�u]ۺ���Np�D�'�Gv�gx*�>�)��`���ł�6�[$5;wCO�~3�N�j�\_����/��������x���p�Avؐvr3?�*��d
-c���۝��-)�1�k�ff�������O�mm���T�0���o|/�����B���ٟfv������8oL�sｵ�{z��ӕ�Q@�\*�Z�Y���Vy���*LėY�� �)�i��b2���fןN�.�M��K��������]W��#& "|���ֳ�e�|��gɠZ�J��@����)�xU�KD��{(�n<�	�\=�s(2~ w>8r�W"�Lcδ����\���'zh H���e��)1�}]֥�L��v� $��F;�E#
�R�i���N�/�Woj�N��3�&1�|�#4P5G�(h&>����L��Q�G� ,�#5F���I{�~a`���kT�;(�{����H�8޶��ٝ�X���n��c�l�: ����Xe.E�ZkHt>�ono?��3"Z�u���V$��)�ߣ�����tzxx033��ѢfQ��݋��`��B�ѯN���w4N�!�^��vW#/�DS
yW�R�!���O�VJ�����w:���w�4�Z���?�x��"�"�[Y�U�`�����< �R׶:b���z��4M��\.��97�{����t�.�49�43{j��x�{��ѩ��rٵ���"Q�xx��y������z�\.j��~s���-H�iM�	 �N�'<���>j��?��k�����́ ��*֙�k�D�cL٧��>��~8�=�m�D��qq<��a��	�3(�NpՅ
L��������;�\x�\c�P��PWA��z��4�z�ٺ.>�J�m]��Kc�H��1������M���r���Y���;{b���L�~��?�;��?њ��h��O����Y�]5 	������A���?�$�l��w�3�:�/D �����,>��w#�g�8;J���B,K��E��"�4DI���v��\#�Y����̈�d��L�#YLj���P~s���{4Y���@3C��R2��r�S��\k%���Yg��`{�p	uu@�q��@u�c�UdDb��X&o��4_Xj����p`��B��=�ˈ3��W3� je0��M�L��v�,���|�����4�� �A���]�<� BT��;ّJWϩ�ךG{�0=�=��i�U]7�I_z4#54�������dL��x<zP�!W�:���)� ����a�SS�3ٙ ��2&I�B�&*��YH���w\/����9���˷���[���z�����E�2D�fZG1�'��W5�4"�o�ӛF�G� o�a�y��?{v>�ܫ a�J-emk�i,�	q&��[W�j���i�퓭�A�9D}T���D=�+<(���1�VI���w�3��jE�s;301���������|���ߪ�?���?|���o��7�^�x8������ً�E����gϗ����O*��W_��~�; ��o���?�8����7"��􏏏�_���/����wo�}�������?���������_}�����{<��|���r���y�cZ�me��X	#�u�:���^׭cx~<=����3�j뽋wDD��r�1�V%�b�j&�C8�] .4M��ý)f�D��r���������\�.祠O:���x������ւfH*�R�a��Cf�*��"S$��+��@NBوG��FU�6�0T�:�~�>�	�\IE͕�]�xo*�)j��aݻ����zy��-�ږ�r1Ւm�P��+�>�7��wW����j�7���zn�on�|��G���X}����'x��|(�m�vE�죈�+l_�?�'�bv��������[�%8TU��bq*U��c��:�p���ө�y�1������������ADL����h�7`YA�Yz�����Ҭ�F�g_[/����i��z&�G��1#�)����-�81J����0�6��7���>�bc�,+|AęTK)��T�����"�F����v�=^���� ���g�QD� �V�T�{U��6���j��6�%��6 ���k>������<#�ƆE4��]:� �Eo]�w���&J�����g/��>�{��m��yZ��z'�a�| ������]���e��[�63�>J?�k��y咲�ajR�f^��,V�u���o�R���"h[�����k�������;#�7C��ؽ�S5�W��.�ݢ�ShIʰ��X׽B$� ��R���O^H�hş�����L���Z�f�V�qj�e��_%����i]nY�����KA�!+�W6�V��K��4��;���o���Ǫ\��<�3���/���������.�ri˛wo�:~]���LJ~���Taf�g�����˯�D���Gf~��U��ݻw˲<{��/���矈��/��O��?��?�������-�Zk-�<{�������t:�%OJ�o�2�*f��C�	�0U�⛂ �����;�L�i�OF.�@p��r���zx�u�4w�8>�"�I$���|:����_������$$d,u�"rz|�\j�����-~���)'�����N[�op����E�+c"Hf|��A���{�Z�麶���g4��fT�J1�#�|
�-��4���z@5�ɱE[WB.Y�2.|\هpp��v^�K��%�?���M�a�l(l�e_�Q���T^�GTak.�7ĵ��)E(�	~�3��*����on��o��*���q:v�����ke���������W�j�����3�{yra~fݻ�Zϗs�>'��ޔ���C+�O�{���(R�-F36����١j������<TD�U�a:��q��;���(��]P��k�"�eξi������N��PCx�-��h�R ���:����W�%�}���p�%f3d�6"�?�܎��3���!I��`FL�hj⓻`�D�-pp��n�(D��
 �e�nN,�31�_w{ ��/�^v�k�����S�!F˄�Z��`�.jH J18Q]|��u]Wϼ�n�l�a�JcA4�u���a��8�ߙ��5��O��������׵Y��[B�ܷ˟�n1
�u�B���ly�O�&������8��bo2B�i^�)��aA *4M����H?�Γ��|���������͍�6ĬOխ���]]N�?�sڀ�ǟ������?|_8C�>�
�psX����? ����۷ok�� �P� ��=|�������&���~Wjy||<�N�����Ck�������8�.��o^�9=�n�7?����/��rY���?��'ʹ�~���GZ1�2�4���Bu2:�0�8�p��!��t{k��x6�|c���<������ ������T���a�����eD���Z'^�����p�Ax��=b]��o�?�l.E�:jɝ��88��ޤ&R�F[a����ƔMd���D�l�(BDDō�&����/���L߾{������eY�j��v����� �BD�[��㑘�Z��I��`e��hב��0�D�(��O��/��x��߸��{����m3�>��鞮���:�TL�
`N�O�vU���:�����m�Ux��G񉲹��BY�Cn��;����A��&��-���a]WN�nd��kX��ֆ�_盙*.��uYE���y�:�#�׻s����ȓ3l9����hH�2%��`�Qb��t0��?���Z bzhD1����H�LmYV�G�P��2��dh.�g��4g�*F��x'�j��f ���L�?ݏr-|�q6�����������ʬ�#B�����Pt�(E
�7�G+����8�l��~9�e���p"�����|�"b)�p�����)�X��1���Xk�J����]u�k���Z���L�$��z`?8x�- "����# ���۟l�T/�OG僂�w�ݓ�|�^�Dc�����E�٩A�͑\�j؁���w{�;o f���������QTDu������߿{���7_����~��I�X5.e������9��no���r9�N�˺���qW;п�!tР���B���3����1f^�ךK��B ��Jn�޻�1B�jbj:�3L�{_���V�«�~���Fo���{Gr>Hm������E3����ӛ7o޾}�$"��ɍ�җl��R�'�|�2f �]Ռ]�$�;F�yi�x��Lj�63�T'$�f\��l:�633��Áe���u7G�j����T�+<��*z6��Y,���:&o��<�t�%���0T�A��+ѡ��)�� y��̀>9��}�#�w����P>`��g�_E�B�պ�P%b&�N^3[׶\.���p8
K(�R�ԔT��ˤ�rss{>����D�Ku8^*o �r���r��� mr��X�\���� �(���a���H6A���t������Xd(���ڼlR�N?��^�"�X�E�@Bn>5L=l������z�n��=�7㗮;����������GVG��@ct)��t!3b63/|��Ԛ����Tx��`�ݺ�WN�|:��e��^����[j����39�70
̞��'��Fϋ���ǜ��y��{�w���S!�L����+|��onfi�BI�z-)*J[��2Q)zW"p.�K����v��V}�" x����6�n[��T��,,�؎��x띸x�>
`��5��)��SC��7�zk�Oo߼]/���=1#@�b��:j\rj�X����л,��㙨���ڊ�d�"����Kc��۝x��y=,��}��������n�ml����k(z��O,n�c���t#ٞ��J�Q��f@������6�>d?�/�Kd �}�����C�����˻�2���b[yU�����5ھ�8M����rY����qY.^L�PIz&�Å��Qk������8O�����wo!� ���Wp����tB��8 3U�*��QJ%,\�t�}CO�nJ��RU��c}s6��ߢF��?梧USԊ��몢1�BN��\���
�5�����(���W�ʧ�C���լ��ꙚŻ~�ٻ�����+a���0s)���:��Rz��ƟI���T�D��-{�g
����)����& "릦����8��"Q��1mjP�*MSE�b&��ؤ�t�m�Tm7�oC;�쾛V��y����vd�E�i{p�m��D��r���&p�A��U�HM��p8������yt��S`��ֶ"`�}]	�Z{�޿����kr_n���̻)ļr+{|�:C�m׍EOVj��c����=U|��V$��>,���e7�
�yr|�@��4�G۞��kQ{B��'O��������Fb$]���q�j뭋 �2u�Ԭ���`d��*3@�5MS��Ԙv��ba��!C{����f3{��7}�20r��	#���LH�Z�Y��9�B��+cbJ5P��e޼!)� OE�c�HC�HUE:�D�Rj-	(K�
�>�� Ĭu� rp�qƈ��,�o D:��R�	�IbfV2҈kWc�����7]~�t�*f\������Ǜ[|�n�ͅ���C��뵐9ac���D�-��(3�i[�'b����њHl]��<�SZ����xq����qYn�y]�f]m�xtT����O,j�<�ۏ� �K���o��Q�*���A�
B30�R<q?.l�Gݽ���Q3��"���/��KuG���)�+	e��-'�d1e� f���#k�i��0 �Z~����Bng �p��#��@P}`)��=*C�u�Ff|��ٯ~������5Dt��r�BI:��|��W���/?����"�z�������'�� �Q$M����ѱ��DR1r8���j��"@p�^wf �y����mU>�z3��e�&�Q��y$����e�н�NVa�Z����]���R��1SQ1���������ba��D��?�qIdfc�����|N���:U���*@���؅3]<k�������ƈ�C��:`������tk� �5�f<�M�]E� ���'�M�5t��YJ^
 � ���uf��y�8�D�!;6���̮�H� [�I&���ղ��LM���3��l�eǩua���g��rYΧs��b����>܆�)���ڌ�� �R��Y��g���������͛��Ƕ�Xv#��Ϳ�e|0�"8�n3D��C�q6��` 63@U��@M��W�� g7x��{�6�PN��lbʀ���c���D	�{�d1��_E��Gߛڕ�J�� �p�優f��� ��I{�/�ı�`��	��U?1B|W���C��4q1"\ϭ�V��GƐtD\^��x�f�QA�����������ݗ>���v�خm�S}��.ˢ*��D���v�`ŵŰ4UEU��p���1Q5<e�z�mtA5�e�F0/��7��@�<�<>�V��SAB��~���?ł�$j�XK51%ĩ�]�b���_)�}�U�>�R�$���,�
�l3���("�n���߽����o޾Y�,T(w��ޜ�FR"0d��%f& �[DZhhH(��߿G���<M���f�|:?�y3Sgy|X�H1�DL�2�=<�g�u��ާyZ��+!��0��-���!Q��M&	������DW+ "ϛ���"� L�u�OV��wU颐5>
<��d3RUf��� ]w���� ��)�s�G^#@��t���0���ޱێ��˼��H3 (T�t�� �.F����EnG�� DB��E��_~y��u%Z����>���������NH@�����51�������������˅K���yE�K�n��а����DU��T'5�)a�J�F����FY}�lb��'�YP�96eVs�� �����a��)$DA�����f9o:Hx4�b�a�]����V�'Rk�\-��CJ)��6 ���"��]�����˗/�e��	PZG /x����&���K�"�2n���6@$D���n0L��bR��}T�-��>����`�U��ēeԨ*��-5�D&�{]."�UI���c{�3�N��+��v`�K���K���#��]������0��}w���#��IQp�	����L������������˲<���3`��)��iݣ��>>�~��Ƿo�=<<�X��|bז�G���9 �fE���eW8 �J`� ͠�.�+F ���6G��X
�m�t��׍�Kr>��=�0l�챤Q�D<҆ٛ����{o.d�P<��`�����Q��{13Q$2T�����\K� �-gN"�!����L31���&y����J�.�Zk�].&&
����Lx������]{�#���ۢ�{���c��C ps�����k��_�~��]km�������"u�9D�@$�7s��@��))�@�40�AZ�$Db�:�� �׏��VI�:��6!��b�Y�R�D�	� H�֚����@du�4��v�S%����P)�p7���I����ۙyr�F6o�D����g���?���}�����6�p�Z�X  ]r�(ڂU�r^,8�Dj�5�������.L"r{������;E�޽ו{���)U���������G/�x�������TU��l����$i��}�V]�wZjED�?J�R)� f �h����bfm�BG�G65'����R'�|4�8= DI��5�l��Ԑ��&��K��x�Q�a&��ҤL�.O�{wX����b|N�w���&�0�n�$�e�#����A[�RDDQ3�R�Ћ�dmk��D�iZ������`��!��[w��`��ο���O?�Tk=��L��>Y���$���Mp�<͓�Zq	��i��+�E\shw��Cs�s)w#[Q|�O
��F!�u Q���=�WG"�����0�B-k����w0p	�2�LfFL�$*�wgG\�'�ʫ�/�i��!g1�oԍ��O��xIS���󡔢j�˥�~<�i�mU��Ee���%y4g�DDz����gϞ���&���q���e%ffF ��U������T�����u)m]ono���+1#2�J�y7�p�3sI�^!�?��iu���FX�'_7&���tC`�р�e"t���Ĺ��zo惩rF3"f/O6z�/��&]Dd�f#{��͛�oT��JD��Z+ ��'1��z��͏?�آ�����a��$b��۶0�,Sc��-[�q����H���/�	m��[�����w)�m�[J�s�1��l��$���K���O&�3- �4*�����.��g�Ht�S,m8��wK���)�"!dQ8 8��mvޯ"�_܀ j73% �*�@fF��D��g����	�].������{@:�{���xs<�.(�.������r��߿���rY"	� �Q���5Dۢ�B���|F���_~��7�|�����?�a]Vb��1�_�U�06�?ʴ�9�vC��ʪ��8}0MTKa��۲�Y���� D@���cI�8e��'�m�8@<cQ*(j�t�,��<BH�v�>>o:�����p"�O�(����pdF"g�%dGb�P��Řg2n+;P�
���r���_��_��_����㧟~����� "�1��d�T1f
BY��)A���(�|�f�,��r1��T�TbƐ�#"������xz|8_.�7��777�/o�7�_�,�S����(�P����L�E��j��:@D�]4r����w������\|�w�S��jY��5^�/��� ������<�ҥ�ֻ/a�bQB.� �zA�6�HF#Sh���{bы������FF�5qokp_����`����I� ��a2-��D_?� I E���+��Ӥ�g53@�����Lͅzk�ԩ�ز���ty��,�[�Q���_������[gFPbrCtxo.�V]|@DUDT �X��Nz_����O��-U@ �̭�d���p���D�Z�*x�9��L����tm���+t��U7e�p��; ����{�<6xa&*L̕U�r���\��BNM{�˥r5��楢˲��><>��q�ɅͬKSğ�٩����	{[/�sk�p8��k>丝}�� 9�+�j;"1c���p,����G-�3"k)���Ҡ��x<N󄙝FW�7%���։Ԍ�j�j�p:]. ]_s�U�t:�� D4�JHH��G��ș���R b4�}x�evW�D4 ��&" km]ׅ#W&�U�D�ijJ-�����]�W��z�\zk"��ݻ���U�XD �k���i:����.�����q�}5WSwNU���o"2��,\�ؒ�+\ez��G�2�"�ǖ0����j�J�$���s)�����KqrcWPf�*�gZPz^��-��u@4���;U	���2A]^#�-侖0]8Q�zJ9�]���������QE$��Tvb6|��/o�H%D3S��L�s���}b���̪�ޒ�Z� �G�N�+'��_�~==L�4�R�"F�c&/9�i��=�# ��0hң��0��!2��Zo��011w�P�ڻv"�����/�?���������w�L�n��taM�8�o����S� �� ��@찇����w�Z�Zk�_w/������~�
E3�h9��Gyx��eY�u]�|>�#����aގ����h�q��'��cT�K�|��i��kڳQ?�1�[�m&��w��6�G� �0���eYJ)o߾���������_�ھ�޻t���kl}��<χ�˅��E$����T `��|�3v>�.����~̐�j-�4;����"���	y9�����C��=��9��U5�t`Hȴ,���k���
fVS�wqV)1*X�ޭ�/��8�R�(Jb�9x�@�og���}L8�%j֛�S&�:i�i�8j�H3�n� 4�P�7;���ѭ�ȅ�i*���vS,^��$+�bίlWQ	��!�����=��;6�a iD���)DvI��BF��NI�ִ�����lh��e���tr�[�;r�kW��o�ff��伾jߎ��j�%�q�2 �D�3]Zo��.MH�BYB�GH3)�NG+r�*10� ץc�<BI�Xm��I�vfr����!��ޥv�B���_�(.������>���z�k[�B��HL��uY��<��S�`��;�I�f�a�,����s)TDEZk����7�aV U]K����oSִ����"a��͛7�JH` �=̶�	#)��޽�N��1<�nU��ljD�����| ���wU�;��u�
�ȟB�o�<%�7�����g���|x�E�c��A1�R�oXi���cng�V��̠�2ֿ�ʅ,p,�w!FGm]Z�@���B� H؈�y��t:�uUw�vǦ�s� pv�hֆ���Di9!"�wҸ�爣 M�;�4������)��b��:%B�|�r�n-���J�n�p{W 0q	q T������d�!"���aˀ��p).�4���ǳH���֙`&�d�Ѡ��k�8���}��KOF!(�h���+#�3M����5t0�k��I��T"��z_W'#�񟬲]�7ꉪ*3 B����LL��BL�+Iʌ��ދ_��J3ׁB�E\s�l��:U����߽������<G�f�S����g�x"�-*sa�P�4��A4UϴB���m�A���L�@vpf���Nd.��F���Z�8?��TM� RA��TST�:	t����U�`Nw��|��k�nZkD��P������?�d\��B�G��K�*�]6ito @E�`��www�����o������p������f� �[�QKnڥS�F8��ֵ��	#@\��Z��n
j&py|W"��D�1zQ�u��s?�Go4����b���%QՈe�� *����J7Äȅ)T�}���Gll���A��3U�R���M��K ǯ����K����[���!�A�"&�9�6:��ٌD�fJ�`8t溈�x�́[&X`\m��a���oe��N�NEq@�[��	1p��F7� @H�ԥ��D���[�L�P�+q�(�2թN��u�QL�
	9�6ʢ���쟍�
��7.�f��Ԁ��?Y��y��TD�������wC��.'a�	��~�F�S�` ��,K���Zm��*B��0J;�yl�9���tw� �*�U�g`{�H��ҝ�q>�N��?P�ECaj�P%Wc�+�"�wCd�����������p�U�A
�ۊq##�_Q��PR�����ų��<�D�؁�R b�z�PLJ��  �?/��s�GʑԴwp�>��7�7��g`�P���d1���m��v�<7t��4U��Hs|�$�}�g�� !v��g�#jTE�k53QA�STq�g��̃��[TID l�i�����P4y7$�׫h�a+�fdqj��3��Y'q}�G�,<�t�c~=���^�U0	bJ�9Q٫DTKu	@0 �vFHLDL�oLޠ͆�Ĭ\2����G�҃PK;���r���XUE�0���|~�
y��d	�\�=��2��ܮ������j�>�޻�&��U���}��t��@p�Y
3�h7S�x�
f���zY���c3�� ̄ �*]��-:��pY��߿���o��R�hm�&����+�l�˺��>u%"gH��R��X�T�y��&���Գ��=�R�yR�g�V������
q��Q^�u�ާ���V�a>��<̀����w���'���wUJȊ�<�LY��4ڈ�l3��K����xs<��GoC@�=gW��;�+Ǽ�#G0���`������|.\�T�C���a5$&d� ���$󽿒2k�m1u�S��e����Xtn �ej늄�t�|'&}�3-��5��3Qw�DD���Ib ��+~�bJݺ�_Ǡp2�������"�ݲ��f":�τąUuY�R)	�Z22sLfu�(���Y�Ot����C�}y'�J�<�~�T�fg�䍏�01\�AܻF��w�5�����j�� A[����� �ܭ"�O�P-�M���vF!"B�7r��>� (iH�LM�{�6:ח��/�9�m�#| L�ϗ��5�<ǪZJA��b(%:H%K9!�1q�S�*'0�J�23�m�_ė&�<+��џ���f�,�ǂ�sN�dd��Z�H.�I	i��D�(�3��Α��N_I�5S%f3y|xl����۶���Z��Y��4E��{k�sCq�
�yd� �[����℘ᑰb����F���X�%��[�Z0@�R0D�-�Z�V�Y��0&b�}G��z�<�wb�1� {W�4���L;?��U�m�|?��� xkIx���<��{Ef�0�!i7 {ѻv`�����H�"h�5w�9(?װ�tFK?����%D/�F.�<��#=���̍l�Qs�c��x'��H4"���O��t�3Sf}ӛs��<DG�&���� �@�ѫu ȥ�̀�Gm>Ow��oȓ�H=Ua�a���QÖdq�؝�ܚz�DG��č�ti��
��P�IA@.ō!Dj�����#���<�000Oy�e��G�pԤ�XdU�18   p��
ę�(�ԩxjl������ �v'�m����ZC]� X��|�����O�������Z�] f�U3 F��%;��/H�ʥ���� S@���������}��?AE��D &6�M�;�۟7�RjT����̧�S����"�����@�"��5�En�D|�r	*����LM�z� �� ��+�CbD`"!R���C��4g��T|�(�Q豙+�5� �b�K���+�L�l"j� O�7P#�0�n���?�f�i�T y��cG[���Iύ���g��+�4�ElVf�W7<eA'�1?�P/�.:��?u������;P`�H0 E�DE\���j}%��Hm��]��-��ԫ<��5Ù%��!��y1�i��|d�p�l��m��F�0 D}/"m��~���d| n(��FL�~K!��@��r�Ѹ� �A%��J�AUG8"iTE5EEL�]���p��Zſ @�}d�b�/��1r
ָ<����B7����%��;�e���k-�4!Rk>�W,@�����0ʦmg�͈ͫYM/��4ϵV�e�LU��G��V̠n�8���+���|��< ��qA�1Z��G��1��:�{�%����6o�Q����[􂰳N�GG�Ƈ�2�s��8��[��4& 0��O�]-ƣ&(X��a�uP�R݅&�"����}Ѹ_?�~TC�#y�a��YN�Œº�Ų%�\D�b�}D\�%�b����[��bE3��&���98����9���Z71Eˌe��lF�"���>6�-����F�;��(;�W޻鈈� �QCE�T��J�Y  Q��"a��
�2lN����5�H�h��O�d�n��lc^��Jf��v���08oj`�����v�cZG/)H6��'�L�E���A�^�y������|'G�s�>Z�������a�~Z5d�y>�u].���|6�"�ޚ����U�Ӌ
(��f�³�#'��v>-&�-����2�i���!���`g����,���99 "�- ��WbM�4Z��f�� ;�� �0�Y�8�h��VP�M�q,���tQ�4%�O�U�	�R�� rjPJ�t3HT+"G�≿4�"�5�\
g����jc����'�\���7�4C�+W=�$���qTX�T=�&Bך�2�z�;LS&h���j�vm���@@d$ء۝D@��b�ѡ��4�~w�W��H�a�k���������go[���'��^�^r�����Γ�ق��Vu��O���G�Q��^�V������"���'�)O��γ���[ �h��o_��A�`;�{OO 
j*]�n�o�R�4O�<*�V�  @2�N��:�D��䬃�TS ���?o"�ѓ'��)`HTEtmMEj�miffhLd����q��C�sr���j�9��~�m�Sy0�y�}D �*�׉b��CA>ɐh��6V�,��rѮ��'���W��-ҝ�l�2ڀZ��ȕ�1�б�'B?<b^�!(� �:��2>qx��z|,��.`��ݽ#��~U��& x#%X�	AiH)BL�����$���O�io�@���q��1��WUJaۛǫ�w ה��6fw��p�a�R��l�ݕ~�/\�+�%���k�m\?�0Ĕ'A"8Y��uO�#$�*ϯ�xΑ�Q��X�'�Hl��Wv{�?�� �Xs�sTX�פ�`+��pUx�u�[�ȣ�4F8�;0~�L��<�T��
SQS�u;e��B�^m��w@DfnTMdTd@ Q��H~xG܀!	���6b"��a���y�����Y��0��&$Ps���:������R� @kk-�j-
T��zYHMx��q�F����G��jG�5 Po�E$�crZ޲#Ps�{ܗLZ�p��~ �L���JHd����`��W��� ���c?"D`KD��߯�d���0�u@�č�!yR.V #�L�l6�>����x�b2F�0�zѰ�nH���HKDI�4�Sh1�(bSܞ�.3��3����5�%������}e|��z��>4N��s����_h��v��z
d���TU1��`��xv�C��zyw!�U�~�)���b�OD��LAf������c/Í���3�a�hA��,{��R�QU?���G4����v,fd�á��z#�� &&�5o��"b3��J)�41�H��,	 �����������a*^��Hh
f�l�����p �g/��Z�|z�6��!P�k�>B�n}�A�����mc]�����
���x�8��> � �O����8�
�b�#�������N�zJȐ�ex�O
�1�#���dh�~�E.���1�>��S�Ts=㳢�5�g?M���!L��q���f�d2�tU�!���7��HH�o]��h�V����KR�o���x�����f -?�LE�#y%e0��13 �Z��@
C�گ0�|�+���8�4u��5�������$w�S��j��\�ր �4���V��t��/7�|�?oܽ8 ��vW�;]w>L��rt���bt��>He�c�v��)��T9��g=�>�x8_-nX����Z��$�]̞�&�!*�uj
\�5����LU��Pj҈ɲº�IA���a><>>���&��OqsKO��^�>k:uMF���1��=B_����sG�D��,�[����g��� ��b�{˃�@'b��T☁#I���x9���PDU�\�p�,~#�a�׫���*x�`0a����y�9 �����&F�ι����	ܣ��Š��ն�<><y: �I�T�η���Q�o#��;Ci0���
 q�;gF����#"!*����������?�o� p�62��!$w��Ko�Z`���(�5��N"�$��J��>z�L"���������y�9�<�x�ʟ>��5nFD���ĥ�l3�X���Zkkk���bEo��b�M�?PŇ�K-\� `��f�d@�\���������ֺ�bj�P��d]l]� �qq�P ���_�����v#��|���>�}���Fe���6�?}b	�?�L�5���`���"]wM`���.f���-Q�G7�%��#o@�Ԛ�	��)���������_�w���F���]��Sy�wD� �шɓ�M�~��o~��R$�l��#M�6�Mv�|�,��`^��5��Y9x
 p������Uc@,�O��L�&�k��WU"CE�t��׏�	K�Ɨ�oTvO!��� o;�ct<T�XU�����k���j�H7Y�������h�_�Ļ�˽0y�H �+"�y��V���C���і�q:�*@ԕy��g2F����[��PS�*�Rk}�����Ͳb��x~\���tTd�=�gq�O�GĠr|V���OJQleHd����e�
�eسg�^�xuz<�?4mV��*h�A1_���3�	��y��ކV��2z�^��[�śC!2�&'�#�?�ap�\,�{��q^a���}�H.��"cw�'_G����F~� aN��?'1��S�xt���������:h!`jw���;�S ��F���~�A�s���Ž ISt9��,�_U�A���E�{�����[UDܬ᮪r+�״�O��oW��u�y��)�O����'6w�Z���ȷy������ňf�5�򞜾�\qB�<y
c�~��uLb��ٳ�>��~���G�Zb��\_3~����. O�WQ�h���g������U�
�:{UeO�53鹿�,�,���ǻ��y�.�%���}����Tonn\�ȕ,K��#����.(�?�{�+�p{���ub�o�������{�s³� 0�]O�O$���R�Y��#��8��7Ll[����<սYvJ��cl�}�y�cA���]`C0$�?�7c��O���5{�x�M�+>�>���q������a�Vq��"%0�4�/ewf@�	9os��x�Y��=��3B�ն� |)�ʔR����B<Խ�&!��~�Z̏Y��TH0�#ӡ��2��܂{3��*��y^o��I��V��^'HL��� ��'��8Tdw�!۔M��Q���R	d�u����j�f������F��3�b��ښ����O�#B���*��`Tj�Dt�\�T �	Ka$B�{���`��
�"D�qA�����L�?HMnonN��*2M��W���ߟ/��Z)�G3c"0�����s�Q�6��<M����qL��`�3��D�@+�1n;E����M����t���ᇔ�f��h���^�����@I�Ň��Ä_���	q��][��(��WV�o<�v���'A�,T���k_u@)���-��=�)��v�`�8at��,�BD3'l���Їr�zO�E��~)L%&�@��"�%g��vK>�%��f�����mK�����5n8�h����O�F53�2p<�*5yR��_�Ce��=���$��l ,�(Q�:ʭv���qa�@ac�F��rs�	���:ޯ\{vn��;���5��y�k��3��Q_�������u�t��׵E����`)Lԭ{y̻w��ي�<4t�j)����\�3#"^d�R�G@lmS�	���c��Thw��������'U\	�*�>�?j|J~�����f��s�[ۍx��A2j2:!��A��"S�.v`�[�q�����%;��Q��I̫B�rw,� H�?���*U���j��ʿ~F��߸�.��;��������4�J�q��� ��V0�B�p����jG���e�d#JtDn�Z��#�K��l ͼT�
f�jf7�CZ�C�%c��g\���!�l,�e��.t��z���I��`�� ��Wl�����A���"�=��/˲�̧� �X�D���ڻ��a)\]�
���^�x��%��E\��M=#�H���Lk-���!D���*`k��(��7����d@XJ��ڛ�("Q=�N���˳�w6�K���:����+#(�k��ET�9����.14���a���E伞[�N�^�\��ׯ}�h���󉔔��N��s��pww7��|>���2�3�;�<6IȈy��E�L$~8���hJ
�%x�:�t�J��asxW;��?�	�B��4���aT�l����	K��9�DX��D�x��y�&�����@l�"�w��'����*��``?�f@�hb�|�흈����K��}�3b�7R��|̸,��k�e�<
 ���e��^��9QeƄ/>�H�,�ZÝ�끥/Z胺M�ϡ�y�!��0�W�M�P]�7�S�a|PZ�[05'�w~�O�/���#�	 u��<����.��+-����ds`O>��XO����4%Trqa[���S���@�x��y> ��|��Q>غ�No��N�7�����ɧ��
t�ۀ�Uf9�� �z'�u]�1�4M�z������Jn%4�G"J�S�5�N˧��E1H�13��!����g�.��3jVS��Oc�B������z.�Ӟ��	"Q����wL!y��bcs���`��x[�83l&�7y���⍽�=&��������t���  �e��nBRy��<��Ĕi����yD2�"6Qק����^�������o	25a�\����0{Gb�N��P�I�N��It�;��.D'u搶��}
$���y�����O��@4�� a�0��R����Oq3}�D��z����W�ΗK[[��VB@.1�b[<4btEAB6�.�(���˗/_��L��UDZk*�Kb���uF� ����cHfN����Q�\�ke�b�@��R���6�|��=�*���0��p	���MT[/s)���	�����tz8��֩�_��뻻��z�\. ���˶���|:?`�Q8���CsĿWsB�_��%G����:I�a��6�uF<9�ӯ@���D|��XmH��sgyM}�	�ݗl�-q�n���@5��0��[<PZ�o���B�M�j��q{�
��\$863T�t  ��F��π�O�w�d ȡd��O! �Zƍl�tw;;���>|����Vfx���q؁�	EjJ~��.ٶ%�.�?R%���.f���Q�}��ZJ�^{^���N�_��Az�WR�R-�DC�W�k5ߪ6TH�HA����2�]9��k���x�|�D��D�7�y�����������&2œ�n ��Bu���Pq��>c�|��� QS����g�i�����yZk��`<�*{BD�����ٳR�g�������, \ڪg�����.�t@@1T/�J��Ne��� �dao�����9>�pl�.��E�XJf��V��ax����.'*Y�����I���v�] ��J)��F��@���'����w� Q�E8�Z̼NO����fA�����b"N �5����3Vt��"@L��{���$��n�Ǎ!p��64�Pc\��3]e� ���i� }Uw�� "��������@�~ ��_����D��&�$��Xw�v��GZ�!�T���+Ł}�|�}I��w��ye������W���爉��y{LQvC+&Åy0���-�]����`���R��<�y>��>������)8��CC��bV�YU���x�ŗ_?�{��Ff���,��<�4�www���f6�jF|�D�!hÌ�s�J�����-�w�"1�4x�����M{�F|%x��ޅ�&��U��uY/�˥��L�������jT����_������_�����D_�z�&���?].'f"f���)��^��������ps{���{����|��]�.���|s����w��lad�1#Tx�K' bħ�+�w�޳w�;����� �y2@6�S,F���ݍ� 59,��zz� ���tu�c��:��]75Yyy�"DΖ���xu����^-(t5�=�$,\c��1�7n0y5�N�)\J�?1�@@V�����>Im����=`n�&*�@N;Ĕ����������wN~�ಎѫc�]���h.08�"���U���\���d����;~��s�ʊڸ�X,W���ƞHfe�h޾{������TD��2�� ���za!.�DOJ*�g�-����5�\��zss;f��\έ��I���=U}|<={�����rY{�Ѳ� �b������o35E�.�D>�w]W�^.'t�B%m�v��I�Ī����޽S�r�}����]���aL�9�W��i;D0��5s���C����%�/j�R\c؉���@rfP��M5X'ˈ8v�Q��Pڨ�˶�@O�
EQ�1��xj�aED�FE�����5U(e���O��`9S۹���T�2>d(�������V$礊)�H	��L�,�!p�M h�C��U`��ע�XU}�{lB3�y�	(\u<��#�`> 6+v�S�(���.,�.�K�	Q�}�loFc1�z%�� @���W��5���~�g�� �PDƁow�^k������BL�����mԳ��AvX���礋<�N�e���uPU�m��4u���%:�O���Ms������?���� �u5S jm=�/�za�����.�wf���pss�{zW"d�y�k��5 2�ZļCCS@R����
6��{��Z���|)����L¦���[�DN��u]�ޗ��mu,�Z�Bm]���|�����+� �i����{_����C[הz$�In�(�FO��R�4��,��6Ms�6���u�pe�����@�h��G pP?8�5=��U���%����M��z�O�̠��e �mU���ƍ3�'��v5�y(�Ŏ`��8\z~dV�{�d��r��R?�5��mz��SG���26hB�8�q�		��e��Z+�q�R 3�j��!�����n�p8�Q��a 	i�@0�0{��ƽ{�
 �S�T�l�� (���:�{vU �lveB��G7�Z]�#W2bS��QΥ�� Հ�����_s�Q�l��L���1ǽ\����e�!p����s  Q}<�N��?)��x�b"s2������Z ]�z��P`+�c��Wfo_D�r8�� >�O�&m��`���.���[�7�c)e�V�O. �}^ew�"F!h�HFD���"��zkޯ�A�%�����P)e]�Ef�(O�����(�F4�G2^����"Jغ!��R��r>j��\��,4��DFZD,��3�8Gf.��-���~�0�<�����%gz�H<�ojP��o`u���ǫ��'�uP�`�o���[�Qxp�`݇�W�a$M�:c��M��7n�i`h3��m���@1� ����w@4 ,��bv�K�d��)�`e���n��W�� ,��̰x0g�t�*:�f.�@�^j@��j�	s������t� �hӞ���_��a*����Z��X�_:�u��!Y��D$�~4��"��N��'��������U,60F�ldͺ� ��߃�&�s"�Ë��={���3Q��N��7o�<<<X-Ջ,�u9��i6����,�<χ��p�J���^7m��ջ� � ��'A�|����+X�Rb�ц`�ϭ���Lː?&���\�R�����ޟN���iYCX{W�RK[ET�i�g����wwǯ����۷��.D������ǟ���ݻ����M���5�^1䪺\.��{������S-�D#��n��e(� @��l�TnIs��5�����dD�Y+ R�#@����e�j��/�+ *�̅!���a �x���ޢee���D!FT����O�C��1��yl�o�[Ð+�>��#�����ޯ��j�L�8�W���*:(̑�T��<��<I`G���Uu�������]`��'P�8���,�r�����kԞ7屳9*Pq�� �@$�ۮ�&Y��HA[v~����`+z�k֮���0�\{ץ# HW$*�X�R�t��ĉ3B�ͫj (��_�������)�8�.$������'��vY$ $*������P�� f &���dfk[=�ݵ#D��\YD��4M�a:��jrYΦv�n�i*�}*��`�Kkk�߽���y��тH�Lk_q0T�mQfmJ��o0SJ�D�\��E���-V	���j%V5�<��g�Tvc�'sT7����_�C�`��1��
1��n d����	���c]��C:�t��	�X:.�|��Ff@>zB�$%�9�j�d6����1� �,�D�W�Dc��Z3cb�y6�1}jfD�����̀����>3� �i�6r�Q���{��W��c���O�Y�����R!@a��o@VЎ{ٟ.�. ��s�vj8��͜�� z_���2hv$��	G���<y�x8�����ndE4�K�	}fr@v��i�����PJ�\Q�@s�1��}�WoBZiL��<�2PQf�6����:�y$�@̋^؋ 1�7���R`b���X���V��s>v>�}�J��DL��|��trL�>uֶ"�1��g�}����7w�|Y[�¡�Ȳ,�ˉ�����Ճ��d���p9����|֞H��*n��z�f��	�q=m]J�`Y�a�j\�O�x�;SsTk�ҥ�G�Zkk_.����{SU"��,m鲊*�4M��.�O?{�_��:Mo߼��S9̵03�ۛgo޼y||\�E0&�"��J��a#���Y�����Y�DD��[:��:�D�Æ����鮸c�k�	��y�U��� �"W[���PF@�����4��;�X�36�����Y�C����(���i���y���fˡ�;[��k���u��^�8ޏcI�C��:���~�5���j��*��n�i���J�2�f��z<]�4��L�@�V(ɆA� `)�Ū,[7��eY}�˙.43D#��U:��7�Z�]oP�C
C�dΝ����>
���1����T���jN	�'��a�Cܦ��4�8�#�(��b�n���� hb� �������b�����9�9���][OV|J��3�O8�+�'���g*7�k14*����'�:�c`b��"&�'��=D4թvA�������xs��"�bj��k��zo뺞�����R���tti"�f�܇��X�yy[.������^E�\QUJ��L1�����S)b���о��̈�����ƥ��̽S)�H�&�wO�#y}���2�'5�X��F�R�9ϵ�.����:cF�F̀d"FCۉ���`�Ú���8�F�Orl P�شKX{^jQS1(�2Q���=VO���aeZl5�
u���ZX�*��2f��-��x'��OW?ITD��?1">}�`����t���8DX�el��Y����50Ba'6��u"@�R'��Qፒ0?�DT��c�Q�b
w^��Q43"C#�܇EA	0�[� #{���{�j�a�H�8}OE}ΉŸ`db��\o�(�5-T0#�����"(z^���K<�P�V���f�Qc\)�5D��y>���O9��wlX��/$O�#��>�Rj��no�?ys���&�H���T��yY�u]�Z�9##һ�P)�޼����r�s����Ԫ���zUe�Z���/��s�f(=f{�w��3!�i���H���4�R��@\����������h�R��tyd����������������~YA��x�T�n���˷o޽~����Co��Pܲf0�Q��nK)f*�
PJ%�Ib*�@Qi�Dר9A�d����9'�����0��#�X��8g�_l�q[�� ��f�4��;L�k�&U�&,�� ��vQ (���z$̬. @k��OmX��HS�
��������e1"��1ڈ��
":��;�@��c!O�D�U�g��!֩�Y�"�Z6�Dh�^���>���N`������.�9�	���m�[�`v#��B�V�1���x���6� ���H�� a�a�H("j݇��_����m���X��љ�k�F�0��1��-��u���;e�}W!b3[��h�R�iU�iD�޹D���|��b�W��Nc'!���Me�VRC�דw�� `䚚���I.��m�'�����X1ǔ���̷��u�{o��.JD�t�����60��<�Tk)��4�N���P���
(������4���S�f�5�̩�:Џ�Ȏ��w��O	F8{�8̛w� �V%��.�䮱G�e\��A��$�x�� ��}��0Q7�Ddl��Dd��i3г��- ��C" �y.�E͘K�|@�����-��.*fڻ�Z��=8	�4�� ׵�)��`0���	J��4�Dq;�P�.�Ư5�W`�v�1G5Ѽ��ke�y���=/�P���s D~g^(�,�_8��E���1�Ze����C�el1��`�4��`�w����n4 B����%N���tUe.^B���C�h'��������1G����!-\UE�YUcޞ��@� ��#q%Z3S��LẁJ��Z�+$&B�.��Fn�c`f2#@C�R|�kfV15!f'hӏD��C32"꽫)!�R�I��/��������/^2�g��:���w뭫,\��"�a���z��9�s��)\�����uޭ>������kkBT��j������ZJav�s_?ϳ6].�D���D���E|ʎ"C��*�)B��&��<��	���(M�T˔dx)\*�����`�b�<����������t>���p8|�ŗ_~�|��w���������x�w>��y�����ٳ�^}�����tRU�.&�%�\
�9�Y��7�<����yBq�����&������PP�C�˂�%�� ��v�螕\}��,�N���3.4�ɷT��Ƕȴ�;(���x�7�d� VJu�%/�,:y��l���٩�I(�zX�d�R"љ�;L�����i�+�V�����ꥅ5f�R���d���t��vn�cPu�f��0�D��-=����-��N��|gf`��d�.��kq�Ʀ����^�6a
�'M$�~�#"�ܢ���5Qͷ�\h�����������wUCr:�e���]`���9���cC�0L�8���П�DW�Q��<��ę`�)��<<�^���hf=�{5	���(����AB�r������x����.����y.)���{;ȼ�S��{����D�һ�iB��:��iZ6T/c ��i�ꛓ��yY�nO�I0�֚�dϺ�Ѡ�M��:����%��b�v@�]~��K��^��s��.�dY@b` JZ��Xy(1�z`���D�
��ő��*s%
��Z����<xD4DRV7���H�,������jj�X)�2zk;O�DW�[�q܉kA"�b�\��� ���#�!F���V~��<��In4�j*ڍfA0���2 ~���Л_
x���HmE�?�-F1���u�Ä�B����C�{2�p-P�݋C��v�\�%����rf��o�^J�hq�T�]�ژ�΅1����JNl Fb*��q�=7����,�+�	&"�b`D�\�����F�0�Ċ�Y�U&�	�­5i�+�=bP0*���ꎒ�THp��к b)\�4M�h�[jd34��!xw��^E��͍����A���Rk53�ZJ�jU��6uf�t���ﾻ\._~��W_}~s<��/H��Ool����ݳz�n��e�����(b���ݠ���<�����,g����$� ��5~�{��x�bbD�=� ����Q�VU���4M�4����Ye.e*̵V�&T	��ۻ/>��7�����/?��h���~�ͷ������?������g��?��?��o���_~����T{_*��^}~w���扭�F���};AxS1U"�j5��۲\,�lj��"@u���B�(���R�_�o��ݩ�%�nyy����#���hCo;��R4���.�{�4���tSs�z㢵TUuɍ���kt���!����k����@43i���x��a�ݝ��ɦE��]U�fg0E2���L�����������h��RDD��1� ��>k m*<J:	��<�0���{��M:�"��T�♌T�X o������ ��.  �T-U����qѨ�$͞[τ���$	�/E�+
�Ǖ�q|���9Ld	��2m��()r�޺Z�O�P�$>:�lja�"*"����T�*�Vߔ;�F����6&C��E�(:�Ə�./ޟzP�l0CH��N�E����]Ln Os�)��}�l];���)g[�����į�6���Z�\�D��ײ,���N���{����W'���hDH�u�`�ƫ뿺L�/�$L㭠�|Y���Dv��Q茙s��#��/t����7ڋF�#�gU��B���=n�9�p�`���^��"�kӒ�o�zɁ��j!:~\��@ �8��T��&DPo��t�0*� ��N`{�5@�qZlu5DR7}hA�"1k�P<c] �F�n�b������a�oS�a"�sK�a9�젏儬�t���e���S�;J�H� D��)��]��8�sF*�Ȅ(����C�M=��ȀTDĸ:	ĄXFo��9�t��B�hҶS!��~v�󦽠A�{P��(�:�PTk�"ҙ�k/T ��L����n]�zs�2��KGT�z8Lf�M:��s4~�!e���U5�烯���ae����� ��r�\~�������������ٳ�ۻ�R��ֶ޾z����iB �v{{���]�[i�2͇�[��9�?���w�^�)�b��u[h�hj��f�S���.͛* "x�*H�SLP��ūW_|���ݳУ0��C ���93ѐ�������RK���٫W�no���������{�˻���_��?��?��t:�y�Z�
�"��������8S�H�4�������݀2q[WQ-��i*ӌ��'1:j#���l�M<����n�� ���[[[[�c�L��hh��,8d��i����V� &�E��ș'��NS��� ���3���y�\f�7���'��4N�E���Ϳ��i�%O��D���*Vm����}�hZh��UAG�`�_�Ȝb$b���@$j-�{TUQ��f3"�����y�½K���+&Vf�.BL(�N�I���&!ܹa  �ȄH����ZE'��.��b!�b.]��!���q��� M�u�8�x�E6�E$�Е�%z|��� �+�!�� �hr�PU����H�7�D P�.=�����ID$U�2��W�n���}��&:r�k�*�ab3O�"�h#�a�6����p%��^���̴N��x0��ri�����D1��Q�x0s���,S��<;5.�6 S2%��&�|:�b!�zJ��F3����zY��A#�x���0(�� UE����_���Rr2g�GB�@ݾ��F�4m�y�*xo�[>$5s��DcD�h}���J� Fl!�|(QF�bՐӺ�qf XkM7����5��Zr�娦d��f�]0�9Usl|�n�w~M�i�$ ��B��hH�L��Z���
^Hɟ1�,0f�)٠��T� F� A�P9ٝ)�C�����ERO���>c��Ȕ��p0���v���ʞ�w���)dD�m �LN8�(� �hw-�X
��DEwE�qxG�ת�HD�c-�b�=��HS�����Bo�E"V����"��ꈡ�ZD6��i*�f���W�˾����P�yb��A��K�gՐ�uz�B��*��v�9c$A�x5<�2MS=o߾��������eYڅ߽{Ì"�����p����v�j�Ì&S��O�͑�<MS���z;_�rY���|���Z*������05�`�<� `XT!BJ$�2�a�p���t8����o�����g���ꀉ�.ˢ�LX
��"]�y>����F�o�4�Z�r~�����}��7�ႇC9_��7}���/��������_���e�����!5Jc�% D�2��X��Z���H_���4M���]iME��D^S�[�\.�_Ɖ+�>ͮ��p���8i��̄]��z'҄�x�E.�c���F�^��g%B�S�LCr��m�W>�کĀ�&X�e�3z��n��C$� D:Q��$Q��/���ʹ�� �yJ�#Lomq��%�a(�6p�Y�F� ��A�G�s"��Ѭ���a��ff
e����\�uχ9�� Ų[S����E$P�]�o=55-��	�M�`��!H�ǌbP7�����Zŕ�ͫ���C���ʭw�(��f��9�F�Gk��Ċ�#sw� !��*I�w
�4"�z\�-*��݄&�z�e�":_�0�s�����ܑ� U0O���'E>��'����%1� c��F��� 0����3$Ch�3h��5"����&����\����V���sk�L�I�J������2{]����bU�w)����=2"�W���Y�Q���xp�i��E0K	i��/o��Ü�u(���DD3�7\�i�OE_�W湚����r 63�>"��wE0��&"�T�*pg�<���є��H�'�{[�I>��F��߇y�x�C_� �!u�H�\.D^�>zD�ӗ���M ��lf����.�Ĭ�����z�\.��`%"��H.AEY��>	�[�B��e�l�0n33��%JZ�  ���
m���,��{P@�c��&@LF��
ahG�2�Qb�RK��E��u�����wp�ğ0#F	,0��̥ D&W�8�6"�:����Dz�JoҨ�b�2vRڴS�^n�Dɳ��� 2����%�pqF썌�M��
R�q��w^�-���Luj�Q � rH�@Tt]���4ϐ=�7bĮJ���QԺ����]�L�0i7P��U��T�}���k������������X���T'UY��͛7�^�|y���ۣZ;/'�����L f� �4�J-SE@S�nw����_�w�ǟ�)M��#f��HT�PMۺ�����'�.�Z#*��������ϟ�(���O�$mU�Hܺ���Z*3������@T�*��Z����w�_��Ñ�+�����w�����������������o��t~x<������A}3k��Z�����������|��i�U�(���t9��u=_��̅р��\�aDU��J���VW7�S�-�!��wByOfuI<p�R�<�A �@n�4�Rn.�nK��Ꮺ�H�;ᡪУ򷷆1")}��W�lT_�{��	���0��u�3��p8��k_�<ˌ˲^�L����{o������{�e���S����h@r``�{�{�̃{�����AN�d�c�A�@�i� a���̍�����Hs z�������� bk�r�����yqCi�46�860�{_.��rq()hDٙj``�3�Z|��x�y�8zWQ1�5
���%���`rL����Q������[���������&e(]�L7 �-[V�[��^�s�H��T�Zj�J�"R���g3Y{�,��rQ��\�pa�"*R�Q �$Z5X�����3�2| �1d+�b�e�3T���g�mB\��cd�t ��崬Ͳ�7�w��N��D��m]{�v3b�đ��]�Z)LĥT �2>�L!jj#�T����6�	@ŧa9}U��
 q�ԋ�!qw�����+31ϼ�T�C� �eY�e�;1�Rx��4MӜ�QE��Ì��̒u"؛+��) q�%"F��V"*�n) �R9����U`���v�ie�7 Ȭ�G�`����]f������"�D�KWs���̒
���p<N�t<�i�������z��׵#W��L"��fQ2��.��  ���߲Aj��d^�� QAs�t����pd{6��Ѿ푧�܅
�:�"\���PJ�*^��g�t0��L�mZB\�̇�N�<�33�<M��8���{o�F�aE�T��R��F;=�_�6��R��J�ҷμm���bB�R[����]+&�j�u�%$$ "R545�>���ū%k�Z�-K���}UUbnmi]��U�{l9HC�=|:=:�*����q�skR
�7D�\.�ZjAd2��I�3:��fj���|��x�����o^����no`YpxWHU����f1&���U��4�1h# XOz~���2�M�+�D �ʬ���ً/�\.�˻w��t�%R.^��PK�n�T ��!g�M�~6ݫt���/>�կ���s�j��D��r�_�1��\	^�w_~��T�U��^?,��:��������1�4b �R�IE���������������7���W_[�� Z��^-�a�[�=�'����4���"�����' xx�<=�Ak���岚�t�n�n�y]W��(�y��Z�����L ]��Y��:]T�Ԣj��6P�]��q�*���5R��0�{\UED$��	S�R���O��ɲS{�'�I���rY.�����<�77�R�4�g�'� ��c{x|X�I���B.�5]����ҥNu���8n"z=y�(`ؚR!@ �5,�(F6M(j�Ԁ%jBD�!����0�W�. qd'þ�^83M���ݝ�����[k벴��`��Z&�Z�=%$G�`���C����.bF!�d��	y��Z�" �R�)!DQw�f�W�:�H�ԄՋUԥ	IIɢ3)!v���:�������u�$��0��uȉ!@�B�,eأ�^ՖeQQgz�:"�V��ϱ1�l���jbk_����c��	��l����Aұ`�.P��L������k�2U�?��.f��&�-"m���ͭ�����"��I��N�~q��_}~{�w���4_.˛w�?�~����?��<\�S1�R)$��3��ܶ��N�~i�(H! �BO�������9&� R����P����#��SЏ..��Z�a��Z���}8!a�y�q]���T�y�}�&�d0W�G`rսx�}͈��D\�7��9H����EW�a�be1dB��X�����0D���u]]Ư�֥��@L[���
����2M�h"�elPJ���k_M�S�f��Hj';k	�	3�;>��%�����V#�W��;B��׻mc�)�@��q�{��͔�D�8�ޛ���tT7/��J�k����<|�(���o���|>��uQ��� `�:M�s�u�f7jv�fk��.R�K���0=��մI��u-���y=o�&CPD��Htn�g��a�F��I�85UUZk"Z�̬�~�����t���T/��{��ܽ�1|�{7D���'����ͳ��77�d��qF @j}Y��������2$@�����|��߼y���������0OuB���lNE �Lxss��ųRk[����r*M��t&��o�n�z>]���~}����q=<��MQA��p�3~���jv��ݲ,f�w���@��D���4M��|>]�
S�ѪH@�����=���o���Ko)/��Y�zyx����򬮿�����o?{uw{w���B}��W��滷���/��
��X�j���o��߿��B�/u2����|��?�k��7D��T�%���vY�h��?��l������ׯ߼y�����ܬ-�e]W{0~���Zk\k)������9����7F�2 ������(X�N�jj1� ���x)��5�� �{7�(ؽ�Ǔ�8(g�XƘF�Ѩ��#r�X13f��gx[[J���֥�4M����4].˲\T����N�U��>G��?��?��ӏ�r^��� R̯RSq�	{���܎�!�m�i'D4R��[�� �����F�+6��d���dW�7<S)��T�r��ٺ,����2�l�����ٳg�<�D���@��cq���e*777�a��ϗ�:�t�s�~/��Y�p!�rss{<�y"f�	@�Y ���[��j��>ފ�eyL4PFgF:	Dt����UU�K���,�@-��/�{f�B�ҝ.h�U�T]��}	1CVOz��׹�`�R����a:����Z�uL�:���U�BO��x%��pK%[f÷�5e�O���9nȄ�Pj��G�)Z�b�����m�_����~��_��9�(rz� ��Ͽ��t�揿�������?�Y�!)x1�$b*v{w����&L�LCN���o���"l���FI���J�w��th��T=�;ϳ׀s!�r�X0��4͇Co͓���-"�|:K�����L\*{������ 8�B=ܢ�t�I�<�S��
\]�����|���,Q�J$�LE�,��Skʹ�����9��B�0��:M�4��<fǔ���Ȗe� �|<�yn�־�h�M�&k��NӐ^�Ȅ .C�1��n���hَ��m�Pj3$w�"��� ʮC+`e��pC��Y/��!73��,]��e���������|8xg�˸���V� �N� Z[���\L�i��E�lfS�UUL{�(�*�D*�*Z*��7�A^U�K����58��D��w�(����غ�)��,�e�Lkr:�;_Χ�c[/]D�#Qkޢ��tk���8�Q�L"����ĢpѮ�!�ޗe5kf���;�Lч���B��zk������_~��tzl]��L9e𼜽��\��x���o_>��߃a!~v�/k��g����������i�B����<�����篿������7�����N�K)/^�x����ׯ%�!ʣl�wO8�.�y��9��p�G�_���W��կ�ǣ�@

.�ǟ~�~}��_����������_���ϏS*������w��������tCb�~<_�z����Yw7�Hbr�\�x80U�һ��j�$��Ӈ�9�<J��˲,�NS-L��������7��33��uZ�:O�t:�O� ��Ŵ��G����EZ\J�MZ���q���Tp9�r��C)x�}3w��Ò�3D1���B[�a�2;e������)l 8���F�S�[z|����x�s%��e�9�mY�����v���ۻi������?k�%I�1]���c���dfeWUW�F���($R�@���O�"|
)�3�d�@w��ꮥ��2+3��-�nf��5󈛙���)������n��z���kd:���u�9���:X�x��>��i��9�����X�����t�]~�e�ה����ح���27�w<����ӛ���-I��ҋ��4�8���!��$b!��<��1"a���z��p��|>�O�Ӻf�=���=}��D�RZ���xcfi s�9��"���]W6�]+l.G�u��>5
�ThǓ\i����=�!�̈�k�T�J�˫��qC��.���T�����$t�k`�)�tK�k^�ܮ��Y]���N�R�k&�/�����:8�y�.��o�_my3���j�!f��K�4M����<���w��yq�G?����U�O���Ͽ��oR��~���W�������~����su����yN���rʹ^}8���k�;W�#���/K?(7�F������@d"⸛v�St|�}'!B�����pa�L�8�FU�9����RJM)i@LH>��!D뺟o}-D �ȭ��F_��rz�ܲ�.���"�U�5/�yYV��W� �Q���4�xs�9Ð��b�W��=�TЦ*1%�`��Z����֪f��v��]*��6륇A���v����⹦"�cĭ�u���j�k��q9�s��S��7�~5�	ko��0�~���c�1�䋯)%/�b�L�)�W1!�Z�K����$�11G�ln��3<��6?vS��m�ny����x��˂`$ץl�o!Q�����Y���T���a]�u��TW�H��8�TU��sx�TGD�q��iܥ�aL��"�)�x� �b� ��R�t�hZ#2��Q?���1'$VSd��D�T��>����>�8�t:��0�&=����;��?�я^�H�n	`=���揾��W?>�������7����j���@cd�annn�?�Rb���ג &��HU��RjV kf& �fD4N�/�a\�y�9���/>_���~��������{#ԇ/>���{$o���ww/��AO���4�V(ZkY�C<�iּC��q�jU	!�6�{h�0kL�-A�:��fԏ��������,�z#b��*k �0ĀK�!P�� }8 �}�L5�<��qv�CJC��94�L���D�`
݄�;> @�Ն% ���QK�����s���]S���U*f���4mݠZ��8�M�F�Jt:��e}~~^�ՙE%���aWJ����8�x��x���������RK�E���е��9�`my�,�Zz�AP�����L��$4췥��ݙ�?l|���B,0���Z���\k�5�ZK�����v��m�D5����'n9�C&G�J1r$dB��f$y3�t>��"���	�6�R���E͙.����*��<�v��֫"�K�	>��¼�� Reo�|8'Dz��]+$,��
k�[7V͑E�7�ۻ�B�١\�j�(���*;e��Wo��R*���;j5w��1�v�I�vNF��bKH��m'�%6MD�/��Ӆ�cJ1%�n=�F�H��z���ӗ����]
��/~�_����O~�w�9����������w?�3)��{x��v2q�
A�!Cָ���}������xW�{:���1�1yS�cN�x��uWՂ�	$�?b !��%8�d1]El����N1G�\���+f���{�)%��L������,z�y�l���j$ �m`��\J)�������ypoX�b���9�����p�sRE��N�� ��}���Ix�"#�dj)�K-"=�S�="6���H+�D�F�t
����tl���"D 2� �T)�<�v�~�q�(�.Uaf�g�Y��x�y�a����p �e-!fZ楔b�H�s�`bJ"�	�ETDF4Uff��S,*��`�5�U�#@-�&t�e+��y�"�F+�*�6�, �.��3#�VR�(0�[d�\r)����T��dp吙5��v��f���D1���qo�C	 :O�-�����5놶
�4 ����0@Ā�U3���B��a�*w\e�����qL�ʀ�xbݧ��������'/��o���_�����a7��4���@���/���d�������K�����l6�1���G===�����E�Y��Y�YA���J���)���B�_޿x��5���� ������o���g���_���O���?�w����ϟߟre<���������x��>�X�u��R������f�O�q`ƉgjV����%�ݰ��e�\�-,EJ�Rʻw�޾{�b112#Gkf�`�mF`����v�d�}kC��\ �����RJ.���|�8����I���',�[����ݱ�5}>�/*�4���Rn��V�\�M�o��9��l��3��D�����۷"�s����4�����4�9���pǁɦqL1�w��y���|�g�ϵJ��L���U�@J�Io����p�λms�Ӆ���� �Jt�,���:�\�;^f��8F������)�8C�cCsnf=�%��(U��>���р1DCU��n��?���|.���y9���XAT��[��y�ɛl)%��kZͨ���w;\
a���2$lñ�^zf�� �%�:f�?�ɢ�Z�ߘ6�5���pHW����o�v��JWw�b��O�D�1F<C)%�Rj)M,��)`���4�)�|dܷ�������ˉ���O*D�"bL)�1k��7	D$z`�����~yƟ���������O���ZP@�c�������?.e���ǯ����ID���e���{o��*�D�-�o��~h���03-%��0�ct	3s�i�"��4U7����2.c߱�~:�KD)�0e�gR��>��c "oeTo�z��[4�vQ/�1���m>P�`��L;���|0;O�<fB��Xv�i^r^��ēfp.�GW��-i���>z�K�0M!D$Tj	�ib��n ���TҎ�(rH�8�ں�˺��ZE��2&o�7�v�� IQ[�)%�u{���ǽzRm-	 �]����i��%��%Л{��u�� �q<�i����4M���'/������$Z@�Z��R +`�(��8��Ժ�˺.�3����6��ֈ��m0�T��V�d���~m�ۜ�V����e�s.9�Rr�RkU��%��(N�34.4�\�a<n�Ǜݴ���Ià�*�!
D���~�(t"�
�2�������D�̥n�ɷ'(��Z�����qp؞��P����?�g����������������1����ǯ_���O��ǿ��������������><J^���B��n�ǻۻ�i.�x߱����� �f�Y�[*8�CU����p�����>�Z�<����f������_��+}��������_�ͻ���\�ZA(���/�����O��z{�������if$������?<�_��ZOc��E@Q�4?\4�=c�tc"��-���xd�"�|>{���Ao�9�JURJ�ݞ����u��x�aC��C�j���*�z^ׅ�R�:�0��|$< i��kQ���^M�!b���[{>�U?�MͲ� s�Thb��9�3Ț�3�;�C̩�Z�:��"@ �Z�Ͻ���Һ���~?���a��%�0N��xx>����k]���a*�ђ��y=VJ���>n`ll2��.q���_�N#�)����dj-�M�\�'�1$��Āh����k7��Ce|ꗪ:⇟ 1��n�`��
A��w�s�ϧS-Uj)1�+��U����丮�8��1!�ft���Z��AlM�&�j���M��yƹ�ۡj>��y6���b4�Z �0���8�0�M��,�"�	��:����۠���jȇJF7��*��Zk)�6ľ~��q�#�_�9e�8/���Mۜ�P� � �0�Cђ���3w��|�����������O��'?]B�IET���-�Ƿ;���)�aM)���j@�N!�1M��<�˲�`��Jm*g�W1m[җ�|Ŕ#��q�
�.8�RS�)!w��{�fns���~7�l���1��b@�`ߪ�}RJ1��H��D��s�UR��0�.X�@ ��Z�4�������j�_5�/N��f��0" rqh�����6�Tk�rk񫙉��w��a�1:Q4���J-*�J�n��)�/�E��o����RJiw<�x>�}tr-E��I}���"��6Ҽ��ΚI�^��7���VZ�LL�1k�T��A��Sr�����]vl&�V��ALq�i���4M����y.��b�W	�;���0R@.� ^���Q1C�º�9��%u����2��jU��m�m��F���
 `cKX�W\�C���AEBbP�sYs^O�'q�a�j ��u�x�*��Y�md.�����~w�����4�4����ݨ���;�����.��5�m��Cu.��~x:��Ӭ���ȉ1���-D��{�����O�ǯ��������?�����z�J�q}�~���wV%����G�����w~��r�
%p��T`���.�0�3�"�y��e�����0��n�1�ƥ���e bC���B0��\�j�u^�,��8������~��?��ե�0�)�!����Ͼ�կ߫�?�W��c=?����!�]!#��qЗ��Y!�D�*�;�[�4���E p(e�����RV�Jɧ�y>/̱VW2Cqw�8���߽}�����U\��b*j��bވ��ND�.�ZkIC�i�b��C��d����B��+k��ݣ����毁h !�`�R)�bSr�j>��cd����Tk����jd�E ̀ 1VE0��漂�u9��x<��Ð�˂����]���|��Rk�*Eq�=ܺ��;�R�w��c�{��r�щ�5A�
����²���9�KgCl�t0��ɹ����8U���]���X �*0!���������0�,��@i���S#<)�T��0�%�ZJ�˲�(���8$�]-��-�j.֞�oڭ� D�܈��~A|��*ޝWP "QPv��8LӄH"E�J�R;��\w�JL�Eڂ~Ek�NȀ�Zm5�c��,B�|2C�)�������c$ �^�{+ّ�~;Zm��00PUB��I�n���Rb�Z�[��K�#ƴ�nn�����/~��<����ul2��|�r ���8�D0�(D뜡6��5���p>ϗ�Н-��F�W-_ �>?�@`�g8`����Ņ1��~�W���֕�
��^�.C }�A�}�^��vp��2�S)%�,��Zj����|�i�v��7*u������M+]�D���]T�E]^3r�	@D�+Ʋ�q�*���xs�FFog�c����p<��8�����2J�����~�#���6Kڙ5�nnn�5�7�R�YM�y;i��MM��&-�X��F@��z  M�ը���f1���;1  ��������j��.ťf�5�0�v�8�i�)���8/��z:�׵8�������	MzQ��d c1Eff.R+s���DEb�fZ�}�����2�B6�V咜m�	�1�����Zj]�e]W�kw����Gm�]�L�������p��77��������ҡа}0��֜M��}�=�]��N2Q55���%��|�M��E�Qp�X�ݴ.��h�/_���>�r��/~����w�ݫOp-�&���ǧ_�����y���w_�|�ű�wgݷT��ĈBQDv����W��Ⱥ. �䟪 ��0���Ev�.6u ����?���<�H�7�c�PĪ��kQHs����/��o�������i8p5Sf�������03o�Cc}���/��ڏ���U����a�|z��@c�i:�T1D4��4N�w�)�qL�Ǜ����/_����۷OO9/"Ƒ�@E��I4�8 ���Z�O'��NCJ�8�v�i������ږ!��M�g�*��*����\�P;I����^��9h��9��T6$)"Zk��y]k-�F�j��*����q��"2"�!�`&�X��_|��z�������������tz�8�:-�y^���/(U�E���v/�T͍f{��/^�u/�]�}��-�C�j��p��qg�J3-"���S����8:K�Ԫ5z��8#2pm�v��4h�Ҷ��-��T��.�� �8è����|��*&����f�n��f��K�1i�aHC���8h�e�J lg��p�4�8l���E�j�3����M������]o"R�u��	 ���
�6��2�.�g[�df��v���LuZ#�ZiH�����ĘR����{���}^�L���`��ɡ
̓�� �i�)Ť�Mi��bcL�$���pLOK)R�p��"�����ޫ�Qdq䠵��j=OK.b��c��M�g �}j�����dq���-���/m c�4n��Da*U�ۚ�շZ�=�Dj6���(�	��&�P-n��c�CK�u]�5��<ϵ�]Jn#"�� �8ppU �]�%11\>\�a'mC��lުq����4ϳ+(Dk�z<�l^�Na�qH��a����j�������f[��\�M)�/�7pz33Sɦ�2iHc����a���j�P� 1� ��[!����Mӽ0'�Klt��f��z��o_֫��3k�b*�j)	�77�0�vSJ��!qH$��k�"�d�4�j����)��!`` 6 h�!��93�4M)�����V|���jŖ|�o噫�65�>�����$s����y^�����E�)����x*W/���8�0i<77��8i"
D�xA�(Kݐշ�/C�͂���5�n&Э�cP�8,s�k�6�EJ.#�1 ��b\�O�^��_���ǇӐv*1O#��������]^�,�~�ys��3rK�#��=o�x�`����5��pȍ��0��J�1�4�9�R��a�ZK�*�������(�OP�nH
VΫi3�6��\-�߽x���~�?z��o�=�p�&0�����ÃTanm5�lD@S)���hN��:�����P�p{{KL!�n7�x��|"� FU
��ëW��_�x������i���� ��ի���<>����7ojWRr�Pj�9��	���h�e]k�9�e��q�43���u�i]��"\�Mu��7OO������L<�HL��a��0)2�"UE�%?����Dnm��"s�J]������O,�\P�N�Ӽ.�����n�u�sd�!�%-��b���Fі6��ͮ���G��hv	��F[+CQ����c�ǪP��J���4# ��yS�9ȡ��-
����{ݏ��7d��b �~�mо�k�1 ���>�G�K�v 5%S��EDJ�eX�ir_��~�!�ۙO͂�|�4#�����I�3���Z�T��b4 U��SJщ(*��:�}a���[rV9hz)�~�����J}D�{� o .S��bL!�\ֲ��h	��|Ts����<ǲ����0k~��E��)nP��N[Pއ�EJ�4�<�����`O嗿����B�nv����~��'/nA�A�Rđ\��<����J�0��tz&Pi3>���ujy�V��-=�u�-�ص��qf"9��U�4�ՆZ~��[���5D��o�R�n�m_�(��!��2�a��*�ֺ�r�EUb 0M#B@D�J�[�cH14�Ȗf5["�*@F��s������I�����,+��f�W͐�bd":�4�w��h5�9�,�Ԁ+����ac�Ȇ ]���Zժ��c�,��]	��(%ڦQ�������&�]4E�TA��-��\� �Z((���2�pط�NL��n7M̼,K�y.��ng	 �tm�����j�M�C��~����o���x���899 �A�U͘��)�*��k�n�Vk3ёҭ@w��cpb�(�9�\�e=�����h�Onjm6v��_9�B�����{qs8�8���l�%S�J����R��`f��s6�ekq �hD�aϧ'3S D~��w2����jy^��T!����psQ����@�!����B`��8�$��cX�B�jb�<y��D!pL�~3Ӑ"�ȗU��h���B�b�٨͟RS5�@1Q�5�i��V��k5DT$�;��1h9$���ho& �a�0"��(`����+��yn���?Aۮf�D|�������?��?��/�����zF�"q$����{/�_�9?���_J�7�ۗ�^��>0�p8���߾{?��RE�*jLm�������ؒ�uY�uM��aL�(\G��N���ڭ���i3�>��R�~	}L3!�<	wg�c\s>=?�\�t]fUE�6���?�bd0ТJ�P����
�(�H-y������R:���q�1�u���'!��ޝ�O�߽EBUadD�Z	�8�b#����q�b����G�b5��P83Qf  ���E�Q#ҐRCH�����̚+�O��.�I����|��9ͬ1U������4M�0����.���6�:Y�EUג�</��n���1ƨ��&*�����z�!�����Tڰ	Co����300bGbR���a�)D�y�Zj�b��Z�aJ��30����Go[�[���W�^�SPE@�;zt�0cJ��RI2���Z|�dO�p{@ϹE7�s�E臎x�H��3�T�=�k�|�������$/��a�������}q�����������_��vӬ������y�"�n����q@��a��� ��TJ٘��!�U;z�|�g�TV�f�~�T�D�(�8M;v.3��^	
6{��?6׭kkf�'y\�[G�{/��ōp"׳�]mZD�\�s��9�U�z�������!���nmி4S"TdC�47�m�b�eY�e^ֵ�CPU�X����Tf��iK��qL�(��iLn$ �s�.�/05��q�-���� �X�E���9C��"��R���H���C�&�&�&�۶�n��Ͳ���gm�iA��6�B�ܗ��������8���~�ۧ�B`z4���tv�RhS	z�ߓK3�ۈ�������C��A�U�Y$���8��c��'HP� ��]`U5hF�N�i�������2A0m����׵���e͋�����,�^�
���G��nwssw���~�w�� ����G�@nG��}j��W�;�>%DE�5��
�~�+�B�jm�t�Fe�2F��� ˲0��jV����O�>�y|*�yf$4&���Ie�������t���"B5qꮩn�'>������¶PT����s��"!��T�ږ�y-�Zv1�c�S�8ć��4g�+�,ߌ��O�>zy#��*��� 5��C�����p{s{<B�@4"����?���/m(_P- ���}�?������W���}����K.R����~7�^�|y���|�����yY��#1�}�^v�i��:��۷o߾������9gu�, �es�� >�a_�,�y9���vi��w	�'������J��Ns�n��ȳ�2i�H���RD�������b��[�}	�}�}�0׭`�Pf
R���m�����̼?�������b>/+0G��ө�J�i�(�λ37>���a�ֺ��/�S��ӊ�e
:Ͳٱn�#�����0���t���.px���eB��9W�=�۵-�����EU�Z5�jj�a8P�QR��e��}<�v���I�)�,3Ⲟ���OLA����;倚_����c�g�ƥPJvV�6;NU�tSJ�0�Q�V)"%�ͷ�72��c�~�EU����?\T�5  �sSG�.V�b�ґF3C��י8u��T�� �Ti�1z�M;Y�A�z���J'�ZS�Sw�1� nˏH��=@0�,�����w�?���0L0����.����t�8%��_?-��{t#�u]T5��1��<?1%��04E���-f#�\�(fVE��8Mj�i�B�,��1��I����yNy��%�n�R�Ӓ��vPk�uA�%w�)}C1�C�ff��R
!,;O�Vq/=7����:�%`Z��81B�)��Tv)�H.e]�<�K����$��Z:��1���0��y�# 4\�eY�u��o�����i�ur}�.�O�Rd��טY���:T9�k)�1��tY�o��9l�ri��H�!�D��=m'�`ֈ�WkIݷADJ.-#a�)�xs<""�����q(�����t���7��� \f5C���М+���%8̄�s.9��b���@P�j�})��D��7�%
��N��@ �R���kf��"�qܮ��֧�"""7����p�v���x{{w���1�*�ְ� կ�� 2S���B�{&hm.�Z�@{N�� �^Ϋ����aG9Wu��FY���40!�Z)�E����xC?���g���;��@�9E�Ʌ��"������󙑐 0��1�u]�6Y"�F�U���x8��Xw���-�Vk�yU@����A���i~^>�ݻi?CT��k��KƲ�#�~|�����~��/������Q���-9oS(Ќ�D�y��������[ى�ļ8�Vv��"��u���_����.�4�#c4�R!���˗�iGD�8�Ȳ,��ׯ_���1���%��aw<:��㴛�����������<�Ū�ЫS501����t�y-u���!�iO��
�؆P_�lD���ٱ�Fe ��W3e"��]�]XgfDmiR���_sKڙ�W,��Z�K��\�l+撗e9�ww�����7%//��6��|>@Ι؅pܡ���sy����#i��LѼ�@�ޭ$��n-�G��=q�!mn�"*�7��716#��@��w�D�J�r,IUĖ*B0#�> �RoE�I�*���=q�	��10�Z�O�|>粺�����cU]�Ej=�OiH��8e)M�j��:"�:w�/��s���r�1�4��01SJ3�ڌ~���&6��:�xt^�e�b����-���p���h�X�2q�!Ę��8�q���^->�PM����H���^zd�fy�U5&�O��KQ��,L�fT�
����o��W?x};���0
��$DL���9s�������}��%TNYAc�c�|>����7�C���
�MP|�� �<LT�a��/�" t�\���[��2\���|��r�{F�ix��4l��-ں�=��������Z��6��n7Lc�uY�e���� j�ZsM)�%B4$c5d$��d��@��D�f��\k�RJ)&5023�Z�9t���S�i����b�L�� �\j��v�n8��kf疖���jk��7n���Z�7�0_۴FK�� Ƹ�홃���aU�55kn/}��$�R��(
�w�����) �Yg滻;bRz��3�RT�������R��1S�[Q��	����#:���b���������	���Dc@��V3sC�RJ�g��]�Z�J�>������A�@�ja��7�Z�T��9��;�zqս�yO:�ǵM ��+
n�8�w�������0)N �}h��]��������R�/G���L�>�W�a�z���݈��ee���4kY7^�6;À,���
�e^��o���׿������~�R�[9ql͑��{q�y�ߏϧ�_���u����
8�sLQl���@VYE�R�
0Q
�0�v�]��X���y]33���׏����7?��?8޿���jyz2����f�S�O^�~��G����1�⋯�z�5NA���PKՒ����ɥ�{���w��(���J���-dF3����o����������%�����n�#��N���'��0��TqI]Υ�|||
!��f8���?===��nx||x~~\�,*�:�Ti��@�j�3����t]��?�03 ��)����@w��FDn>�c��E��˺.���&���L̜b��=`I?�	��T��}�;����"�z���<����|zz|z����ׯo����1����t:��8�eYO���<w�nX��!1z��M�-v3&n�̭a=��.��a�ap�휋'aW8�7�q�k�>���e�N] ��s,�j�	s}(�8~���a�!��1q�Ӽ�J)ym�s A��P���*BH1%v��=���~����j���g!�D))F��Ni�mf*��m*U*"0��K�YuO��6}����o�v������V��tPDT,�����yH�bZ�\D�L4o���o���_hH%���;��s���8s��0cE���_����4��^Cؿا��;o�����^�O�x��߼]1�q*�`���I���9D���1�Z��)|x����|�JV�2e���8������j��J} �+��vآbq/����T���t�>	b�򯞈^�7>W�� w@��?�ZN���8�0��9��A�n���0���@ ۚ�h\K�Zr.kΥ�"�405���{?�ޘ��p������ˑP�J����5���Q���>�� mײuL��j���h	ֶm[����Z 0���`�Fp���x%�N�=݇zv�ҹ���V��~��e�8�4�!Ř�q���0ļ������yV�����k!�D��#;�U�Dᵨ���@��I8J�M�tU��3���q�u<�R�nI!U���Eb��'Mg�yꠊD�k+��q���h�$2h�t�lo��ŏ��j���4�Ӵ;�����n�Um�y-Ej���e�·aK�D��t֦#r�����@烘��s�1}/[GbLC�:hb��1�*�*y-9��T8�/�?����;}�������a��ݻ�yF�����������;<N���������g�S͉�b`�H�S��8qJ��!p�)77Ǜ�Ԇ�]���������"�ꐒ��)M7����'���������G�,��_����S��bz������/�������O������&�U��D���9*f�i���_�x�Bꖥhh�U/�{�����_KzrΟ��h�4~�Q)Uju�(0Ŕ�VU����\�HQEo���\J-��s�W���ӴK1�0�wwww����>=?��`�6��%6S��B
����u�Z�00�f��͐�Lq�F�t��b`f�֘�Hu���!oź��Ü `� �۱}¥�:���'�| o�3W7�:�N"����i��no?z��z�����Ǉ���&���R�|>y���DlEQ���Շq���z�Pb��-.�;(D��:,�Ѥ%���[����%:�޿���k��j�;_�_v��9 �<������0�X��x��x<c�>A��}`߅���&V=��IG�Wp�5�[�?A��"L�� )�x�v��O���V �*`ۨ������tfX{�Q	^4�j�7W��7!��3�����T�ٝn9FB�iC�	r^�y.R<vo��_�z����8Ck���-�Rj��	��y��������||�w�awT��3����o�=��˧�	O��<���4�IL�T0=�����픦�W5s��]o�њ��ap�B������%u��o<6���X���μ1w�j�{Dre����W@����V@�2>>��Հ�b��&�<�Rr^�j5�����@LjNLa3���L���Rj)���*"��?( �! �`4��x3MSG�����W~6�n� 
��������u����wW:���)�P#EE1s��F�q���>@�R�ZV!�c��|l�羮DDB0l3h�n=�n=���ؾ3oo�qdb"<���R��R{>���44o��7��^ֺꤽe�VD��ci3` B�K���vH)��Ա��d�\�g )�F04O.U�k ��Lf����D��N��)�n�xu´��ȸ\"ό���i��4&b�X��gBL��L6V��DD���䎭^E7K(3''X����셋!uZ�b`�ݸC3u�R��`�I6�RmY��y��s@@��|��w�/��������0�_�}��I���������t��q��_|��?���NJMԔ�9����s)5��c�8�9 
���\J��Ϡ'���ǇW���IU\r�a���O���W�������O������������ :���>z��5��������h�B�V�����<�kV�4�a��w�/^������Ӷͩ�}q[�&�֋.��R� N��Z}��L3D����8�˚I[X̄����|:��8M�0N�8.��8��n�9�<<<<��|���X "�����*#�CL�s.���I��=��`nq�>�:��ȼ̵��y�ymB�ٜ���W�0@��m���r�}��@ĭ�I0��p��漬����v�����0��O' L"Xs֨ �iˍ�l�]�\>p{�B�����a�|" �<�ܨ�;?��.��s���e!���^Ԏ �)�ͼ�ww}	�ww3[`]�u��8���~��!���4�9��9�e]j/A@�lͫ\�Z�=ط�*Zj�ܴ1�| 6��0�q��9�uYm;*����Z`n7\��jpu� �����M
jWB�W͠�nM�v9>�1i�x�Q *�&Jf"�U8ƈ�)ƘBL�UJ�~R�j�W��sYTu]�0�n�{>�ל�\��)���QD
�b���������?��ǟ��ُ���iy|��������Χ�����匌�a��]��Uk^s�2�S��9*W��!��G)���@v��R�!qh]oɥxV���E���^�ݷ��jl�����ښ>`���-o��i��y���n����HܓW��r1�q�aH��-�3�R�k����J)�\� RdfCT���h�uc}n�n��a�qLip������oT��_�Y�#BtS�~.\�(l9�y��/��pd������j�rJDi�V��1i��Y�u]���yB�[�*"�5;Z�+�Guw$�fv9$/R��x�Db�1��期Eѯ��JDL\E�v�A۪8g��@m��C�� ��$R�,��g�(�L�秪 h)Yj�����"�d�˲���a ����ʪ�"�fm�w��>�Q�
/7��4�̈́��4��8��>��0WU�P�j! ��!��ʝ��F�1E��/�Pg���:�A��%ž��c���21���l���|:��E}x��Zk	C��K��O�x_�OU���?���nn_Բ��И�a�������������yzQ�����Hà�Uj^�<�E$�6����ͺ���kɹ� )���]xU9������mr[�p|�f����O!���_�����?�����oK��x{��l���������|�H0�pJ�9��<><�}����!MӴ����w��O9&����KPӮu�",^:��0�V4h�&5�{��3^��{�U
���|�������p3�~���~�����|�%�Χ��H���P�J��a��Vfm�B#Q�"Ꟗ���F�c�S
�1oj����,��%w�2�îpȆ¶�{�b�
��b_�s���pk�C��A�T������n�{�������PO�ݲ���s���<�gU��h�����DS�A��f��0�.p0�Z�ϱ�L��]�	�:��-l����;m�Iu�1dSݮ-t�Z���jht���\2{�)x��5�벘�n7Mӄ��4wh3/��Y�d���#���65��~-�����ADC�f����\�����cˌ/'Ƿ�ld�-��O<�k����x�C#jy6�!u�2#��Z��
�R��pB����S4U[�"�8�г}�M� ��"s�%���<�M�0䜉(���8�����V�2/���/����>N j��z^�y�EI)�y]� �i�1�j�K^�J�j2ϳ�NӾ�:�O~uT����D	��w��Ӧ�Q�1"���,� ������M��蚳�ݠ-��
Ş5¶)Z���/���g�#"�dh"f��R�3�x�&�u��b����b�D��jU�6u��B�Ш/�%�4��8��� 
ִb��+����v��r���	��������ҹX�7��[~�tBt�#{����R'�Go��vU���1��`)ًe�&^�9�M��W%k�;���h�x�i�h���{���_;M(��j�����nE����F��7<�����f20���U��`�e�V�:�Щ�g B �˺���qMCSJ����u-%�!�� �xg[�7͵5�(oI_8!��~�SJ�����n�&�CR�HAŊ(n��6�<��@�a�!�2_��"_o���&vH�O�z��-���p�UGbj�����</�Q-R��A�NhF0"�2��������>���?��~����b)9�t>՟��?�˟���|���lzAq'
d"�%���oYV�P���y�"�Hb=2Z�w�|:�{��ŋ����s�}H��/�����_�����O��G?����6�,�׿|�o����x��a�qw�{*1�毾��������!�q���n��혹���O�~ 5���!�[N�E3�eA�n1�x@Ug5�7�G{O��*��IUv�)i��)C���ǧ�'D|~~65 ��uS�ٶ�(�C\T<9	���Tޫj캭B�J�O�Y��$j�Ҙq���ۆ��`���)�><}�Q��V\����>��dKN�g�^�*��[C��Y;���w��������f("*��~'�.��)��V��{Z�~xۈ�Ĝ��� @TJv�Ts5�\t�v�Jڪ�������y
z!� �բB��"r�Z �A�-�t��S�y�G �FD@���N'��0��p�r�&?N�u�]���V�XGn�� �y`t!�M�8:�-"�8�M<��7���_��vS��W���>�/��sWɍg�8
1��˲.���P T��0Kq�1�0�y]ל���ZKug;��)������(�>��se��� �H����l���~�&� ^�%�\UC�
�tzN�Cq�y]���~F@���� �G��ÔK�yE0�P���d!b � l�t��ݯT�����)���t^��B�m�j�lw��x�"��vи�@s�8�7$�7���:�.벮9��>ڱ/���Ɏ~|�!��׸���&/��UDE:@�΍n@����l�L^��[_��[�=�x� J�9�xI�|q^1z�ߴ�N��Ҷ@�*"eY%�PHS��cH)�Ⱥ�e9��� P/O̬�A��3@ �r
1p`�U�@YJ^�eYJ�Ĕb��"0�2ۇ;w�0]6)p�����Xv����&� "lǯ��F����s63-������5��8�����,mzhɹ�\1����Ԝ�N�,�i�����	�̼��������ܗݚ�ڪ�7���ahD膓�H[tRB
`���6���.{��:���@F����{��kKD��n�cL�����lƔ�6�+�+�g�7�����>�����wϿ��ͻSհ��K��80�A��,k~|z*�M���|�W�����}7�|���{DA��}�����+��-r`�`���WO_��7��ſ}y7}��ŘƧ�����73J��_�p�
"5%�*�|:�y��t^�a�M�p8ǝ�*)1�IG��f��X�!;3��j�e��H���n�)qh���h��m��@��`�	K)%���	R��n^�zu8�B�|<ެ����N�S�����DiB�j"�z�� ���B�r,�3�R��tZ��L � ]��>�����zE�p�V�6�k`�����og��1��8��t!~�t;�$ꑦ��J�U7~2[��ݻw�y�����v�z��Z+1-˲�ť�x}p��A�r�rJ�8f?3T�d tL�l��i�a$��Hڕ��]�y�Z�nvhm�������N%�V7�bϕ}�Yw�hɭ��������y.���zc�kn���Zә���t�t�jx�˩xN��Ap������*�[a��O�*ﾊ.�������mi�gf�ߙ]e�h.�135w	"�1��c�1�8�a]�*��뺚A����8��J�9��*��j��3!fS]�o	�3�UoH�;O��j�R�i �u-9�����Z���mlbHb�����a����0���K#��2��R��\J&?��z��`X��@��׋f���1�	}S�55�m'�֨�R��wq�圻�?B��۵�׭���_QT|��V�Zs�r�� �7�b����<���K1k�`f�Z`qhW̜�4u1dǑ)�7G8Eki�<7c��:Ǯ���p��
���m���qc-\�h�e�;�\��9��x��;#;�Ĺ�T��H�%�Й�����S^W�vQ����|����yd�!2���]� �u�9�A4�^�Vf�Ȩ�;�Jkˬ�"���Aӷ�S5�{�p^�"uz���|�.�j�C$� jX����q�ݔ��b�R��eY<����Re�AmsF3+"f���n:����d>�p��}6�qv�/��\�\�6�"��'��e~�6L��?�ܼ�����7%cC�6�z;S�j��/:�FH1�aDv�R��<??=�Χu�OOO1�!�Ӕ|�12����:����I��2��is���Ʊ�r 
FA�ɤUe>��D�G6�����	�B
a)!25q�����������>�9"� �"�q�^��e<��ï�������4��Uq��fw���}5�*R()-�ӛ�o�OO1���������8C������v�:J�/�^���W�� �Ӗ����d�0s'�-�A���������.ղ�J��|��9�v�W�^on��秧' ����쮄�����W dv�>8��BH)���m�cD�eY�y�&ks�u�2z��M��m�uRo0qg\�����6K�귾���O&��z��y�ל�a��v�8�|����CJ�L��YEZ;������f�B)rf6/Kqks�>ٸ��
0�e6��R "HU����kH���Bp�FB�����;r@D����5X@ �Q��ȇ���6��B$f뺆}�'�����U���G��U}�jͻ�;.�!=�# �/v��M�f>^9"A�7�������Vwߕ�֟߅5^��7�e�&��\?�/׵ظ�;�0!��Y����!Ƙ��p����e�q��I��y�ϵ��9�̙|�Θ�9Ġ�h��*��jF���͐x71��cwj*�9��AJ)���qH����ngf%��a��{�7��7�����a��Y��n�e����2f@ی�x�u��K��@K4 1#C�&�ۍ�7k?���ZCDD�Hz��*(��S@K'.Rd��[�|��8L����*��*���2��ꮳ��3�0N�8!��bLX��M���z�@@~A.��u���Z�M�hf��ؿQ�^}/u	��G⩣/
0�3��h-��m�{&��ЫfKw���Y�R����@�y��eYל�j�~��4� Ƹ?�i����B-��RJQS�0����}7z�C��ۭ�Eo��!q�Xw(w�WQ�}D�ȇ���.�vIU��ǖ���ff/3T�TY�Ut�b1��j��,��j�U*2�Cm���D��q�v{�)F p�����X�{�b7i��O����AT#c""���9�f���z�b�_<<�7���P���f�C&`�}� ���qûx:��y}O�K@�
�шm�a�T)E�<��0N���j%�q(Uk�j�����ÚDL)����*D(Z���Zj���d�\��k^߼��������V5XK�	���p����p'*a�D6�D�ј��b@����͛7_�y����W�77��.��r�]ݩ���9ڙ%�@��$m9�ޙ�j�Lz�ˁw�/3SQChC��!C-�E
*��K^���a�;n�i�vo��t�*˲�N���G3����
fQ��CSJ����y!�ZJ��&V������b�gK�+W�k�9_�x)��jP����g9�)�[����߆.)5kԡ����B��~��p<���u��4U��l�� f��i:���;P���u��Y�x^�M�"[S��;Mh�û�+��2 p>k�,̤��W �԰��Br}�5@U�n����?�M� S�
Vk]��V��C��΅ؒG�Z>���JC��1���T�f�'�wƼȽ$o>���v������c�j��ա�-�߶R�B�a��p���i�B�*l"!��A�*�T�1ƀ��>�� [���08� v%��H��/�1;#�~�w�H)�Vi�u����2!�g��R��k�,N�k�?h�r��Ú��(��]Mi��4y�R�ln~���8���U#t]�w�|@T�k��*��W��
3P2�	�%�_P�*�O����-a�g~d��T.���H��YQh�H�4E�q'$x>���ɪ������a]W�4!D�E.��^o.���RҾm[��.����،?\�[BMN��*6�Z���w�_{�Y�����힘������Vi��!��wf�8�.7/���\���B��8NS���譪O�gsR�)m�>�>׻�q4$܌��9�?��M���}U_�����RF/���ۋm����#0Y�zC`"dB5���k^"�сo��b�g<�ggX6��=�C�0�42�0777�8nEQq])]!ח< ��[нW���~��T[~/�h����mu��Q�˔�꺾������+1#b�)Ŕ����q^�Z�����x8P����j�!��>�q3Sƀ! sU3N�t��Ҍ�c!0GU��?m0��:��E��}��Z%�xs�),y	�l�RL4���t�����4FPC1#�� L�,������)2�ݽ�q�KCHָ�>���� �i�5�hd���O8�	�� f�΢K.a������	C-���^wk�n��ֈ!�Z��7_�N�~�?v�����i�k�<M�qk�1EDd`h�D�n������x�1�$���u)y��b>u��Z�2ߢW[پ�)"v�𫥎=�@9o�u�{�B�%����Շo��03r"��YE|t�a�?o���8�i]�̪�R
1��sV3&���nd��MKΧ�,3"&J�P���C�b�V\��!��Ո���Ϳxѵ8gWj'B4 G�8�wT��z��*1C?��s�,0��A�e��� 8�m8=c����MRj�y�+"��q�  �B��Zf��nJ����l��>DP ����Wf�I��=�n�AM���03U�~���R��^���[W4`)`�cB�"b��c�H)�ն��٬9z @��|>�8NDB�Ɠ�.�x��Ch�+D͹��HH�m�{�p�����bJ@$��Rj)��q|����@������ŷ���7�����)�b?��] "��< �,'clo�s��GZ=�(��;,�Q�6XEMT�yBo�̤��B<+��c�9�Li�Z��y]W@p��8�R���'R%�⊽���#!C�M��4N^����b�·c$o?BcK]�v�+u�V{9���WU��*�TU/���׿?�F�U���23��äJU�(R�ݎ�8����4N���.��`�bH��8�)&U)��L��m��+0q`���4�s/�Zl0��7����
�md� �g^�vd����K�d�5����������3��f��"&w�;���4��q���@!�a�����4/K�\� ��:�1��$!�Zk)ݭ�Y�:��(@�o~g���}��w� D1������̓f�������-���@�VǠ������1�x<�q�9���R�Rr.�0$����4  ���)X��TUjQ ���}�9��R�c)9��||&  �Z���d��-Dd�O����?����Nj}z~�12���h�5�
��P�Z���
�R벜������^�F�53P��9��0O�����;� }ؑ"A�JA��(��YL���T'���-k��G[JW���h���f@Ujm#�j)eY?N�8�i������~X��'�:�<�0�a��������9�������i��0���}ҭ޾t$���?nc]b�^��QU���}D��uai�
���Ի��̓�o��9e���}&2�������q��������b�����RK�)���q��2��yYJ-N�x��X�$Ĭ56��m�e�� ���v ��o-�2?\�S안�"�F��5��q���Qɠ��i S��d=}k3g��uf6�eYg��lGBp�B$�<ET���������Q��"��"�D��n�=�����sJU�&�.y�պ�j���w����ݕ��z�|}�����s���v��7�b���T7��R��Ę�qr��m1�R�糪�Z��3�5���3ᚮ��)U��˚�ܚ�ډ`�������1Fs�@*m%��xǭ���P��q�#�*��W*�u�b�H{�b��o���I����8�`m��U����.'���
4?&QaO���k�@H����}Vd[+�"����'{��i�qs�fB�<i+um��Zk�#T��R��v�H���W��0�A�8x�U�Fyg� b'��*��/���� R��"*���6�Q���J0TDl�Xh ����}�PD޿~zf�ݴ�������Xj����jV�8�J���
��6~'���=�Z2���V��H���Z6�c��7I" �msw;��k	/�RD"S�Z��M�����W)���L�D����e�f��u]�ֲf���Y�0��4==?�糉:��g�M�4N��wT5�,��k�'�'	)%&ʥ�(��[��B��B j���?{�*�Djf"9�ڨ����Ʀ�p@�Z�լ�d�Vr�6�ua>b{-�I�
�N�8�aH�r6��9�O���x��n�z�%B$����������q��� "|zzQ TU��,*ZrZ,F����uju���a��O~���o�!�w��W_}=M�W��i$��-�)�f���_��̓J�YU�aH�0���M��V���II��Zf���/�����D����v��4͚���奬���#[N�03cFC�vi�Ւ�Y@�B�������T���� c��0N㈁b��>������t*��������nb$��˺����|~���@a�ߍc"b�_
��lc����Le/,A��}0;�tk���σ-�z������b;�����3�)f��z�ڙsz��^^���EdQU�G���p�R�1Qyz|*��aH� f벜N�ǧ���,"!�qC��}�{F�Zj�i%\rJ��{#V�-��#�� ������W,ym�x�����1r��\m?�Z������:�a˩��Jb. �Ժ�K�k��724ҕ����^��?H1���x�ڒ�^����QQ���0����&��z�4CU���&R<�3��>B�_ժA�������m�'w�& �_3[���Dĵ��?���k��y^�մͩ�Ɨ�Z�<ϪS�Dkv��R�R�Sw�ZKYץ�:���DUA��Ӑ�a:!�����J�����	�)8[�j���Z�W��U�t�����b
[��/ԶC��LT��|�<π�~�e�@K7:�ٲIq�7*~hK��Y�*������w����r�F�Wu��ac��0�(R���`��e^���h�Fn��n�TŚe^��g��uV(!�}�A���Ew�s����q��Y��и�U�Ⱦ\<Pe	��)?Pm��U*愁>w�wo����Z�Zr)P�t9�fp<SJ�x��y.I^���Rrγ���D��!F���=8w�A ��Pͤ\�03񏈀����� �U
�U�cU��"�a.�עS�*[sX#U�Bk���<"y��J��K^�|�v��8��iƔ�4��|>K���a��������\Jq9��������Ny�eYZ׹�&PsE�H��I�kR�J��d���X62�^��?ޘ����oWo]�H QQ1��m7�@1FU(�R ��v���z���C����R���l���D���sy~>�}�6��O���0�_��ホe��b��F-T��!����5�\r�_�x��'���݅~��o���+"�ky����?�XݧW�.��h]�Z*0R�u�粮��ޡ�R���"G�5�9�DL�Uaf�[cq�}ϯ�������}���9d&S]�U�d^�_#������)��*E �N�o1 ]��"w3�i�x6"�M��x��L1�Ҵ߉TbB��q�y��޼y���h�!$���c U�>ŀ�D�o-/y�_n0"cCj�m���9�~iD��b3G��
�2�-����'=�*]2˞;`3��\� QUU/���;����˲0�n�{��;�{zZr������t>��\j�������Pq��v|^F
��Di�+n�"^��b���.�(���m^� }�C�t��i����gf��* �vpDĹ�U�̞D��a7�#!�\�����i�O�Fij�����ZѝMz����p%$w`Q��_�/���98�gȤ]��� [۴c<׹hoH�/�MW� ��Dw�T�>��V��D�N��FG�e����J�D* �Z<�c�KZ=��"�U��"����ND"/��/g���R�9�Y!���zb
]3�L�:�%�I���JDjB̨f*��2  �"[[`�P �!�����ֺ1�Zj}w~�M�ɭ��4�&����[�[7D�/tm�d"�Q��,T7���7~�^S(`{�n�d��9�R�n��i�8���*�kY����e�̶e3M��f<�%&\�c �t�F�w@�n�H̡�g�������h���ސ�2GD/�Q�a�.�׮mE�<�H�"�efD2�1�&R�,�`
E򻇷��|{s���jտ�����ǧ'	Ģ��A��R}��6�&JLL�ƨhX����j�\�3��vd���2���g��(����X�������7���B9m�\���-�@[�ֻ��v��֚��|>Oô����~7NӐR��� 12S-�����0K)�B~*��d]�� * zA�X���=eff^ ��Of�1 �JC����U�ެ�%��X o��������W�Epr�2��0$1�8���*3S�R*3��}VH3~v?�����E�9�s�����t6�eYE��onnno�r�D8�O� �CP"j��*UD�Q��ݔvt����O?������o�˿���~�T��|~|x���>��{�i�U���0��ES�p��Jȥ�Z���GD}8[���J-ZJu>�֪��n+e���f�2j?����y���2�ྐd�>Ђ��j��m�j��ʕ��W������D�&G7��c���)�y>?��Ǉi��������²̻��+2������W_=>>��9J0�A���U�^���ŝ۫���V��<�;?��-�H �ڸ�Ƥr��yCe��^-��5����v�W$۟�6
��4���eۄ4D(�,�z>�����ׯ�c4[�yY�秧��5g%DF�y9{
Ҵ�>����і��`��@��i�5���nW�L�q%Dܚ��VK��5\��˿%V���|��m!�f+ �R���)��V3;!��<�Z׼�N��UQ5�f�
]��Xv�#n��!
�4�R�\c]`���~���忻-���IW����W�`�j�{Zi �wh��K�
zEzCd��C/+�߹.��e�s^Ѓ��#&�q�Ɯ˲��n��!�g��\\�{.�받I��B���>��b&D4���y>ϋ[�T3m�Z�m`�ӰoK��("m`��>��hm�Q��G ���5x֠�n]�x����[��rS.��M�����^]{l�����2�:�m?�����j���\E����2j�����|�� �C�N�U��&MpQ*��@����h/��@�) >���e���;m��x&�vC[@��?�d�RM���NG&�H��L�x���A�`��U��)�K-���>=?��~9�Y����O�R2!{�Fn�!�*(��U�MF1a!a!#4l�)�{y_�^^h�!3;)�L�����N���]�%��-�i�!/O�Ź���AN���b����{�fj@�"���tY�ǧ4�vwww���#���ڼ��OO��[(��-���^3�t�JK��P���^_~�[�Bh��&5��\�+)��=�g�NU��3Q���{�jn�G��AΡT3`>Ak�x�FK��a!pR J)�<���sj��@ĥ����"�p{{c:��%�4�r�@A����V,!�����,�|��n�?Ѻο��/>�B{+*�����e�߽y{<�xN��٧i�����&K5S���/bpS��j#����˂F�T��~�"�B@B�"�b��\R3�i`7ͺ�2�Z(9��ZE ՟�=t!im�R��n,�-:�6���{3̤%[^���\׵�zz>=�w��3/�*R߿{�c��EH�5�z�;0�P�5�B��.!۳,�y�<&��!xk;U��{��l;��]f`VW�{g�N�n�EAfBi6Q��o>)ϧ�;S����l�LD���s>>L����h�����[��/���֣�Y^af��Cp4�����-�j�6hg��9F�F��6S�v���)y"�Ii���<r�J.yYVS��1�Xbx~z~~~�eU��lt/OزF�-Q�׿�h`����-�͝~[O=O�mW��̳x$l������;wQk��j�\����
���E�������	3����v�+�j��M�O��J��Rf��k�ֆ���RU@ѫ%�ɻ�fj��6FeҸ�f�a6������t֫�ۿD����D��-o��Y��Ц%"005ҪZ�r&bd Q�.���0$d@i4k�mFh��6Կ�@�bU��.��.$T!��l)�{8�m��Ҿ$y�$Q�,2q�*����i�������|:={�S�b���&�2 z�G�6�ѿ`�p��9 D��J�5g�V���E���[=� ���E�h��9p�	�G��"k;�T���VH�f�����UP��SeYr)y�&B|~~z||\sv�>p�RU�9`px	}40"��Owe��X$@I{��.~�m! (���s[͆G\Qcԑ�3L�u�o�����|M������	���T���j-�[ϥ6,y�F@���K~>=��'�5�ދG!w�궾�6��iS�#���VǊ���"�Ԍ���R���&f�|��[����b���e�������W��l��G��@U�T0����e{;_`�����c������"�8p�c5��Z���gO7���ҐnoooooK"
\5m!P 
"1{95ëW/k��n1<==|�՗_}�U��3V �)��������8�a�aLX{� T+z�﹋�9��%KU��C��J�N[/���@̈m����1�52;��j������w�3�U�c�������
TG��s�o �$ �g�.�jM�q�o=�ϝ'3+���㓼zT���*�����կ�#���0�L��B�n%�W*R���t�m�]���>�e�]	��t-�\�m��C���ۿÛ[���n�aB[�@D �r�K��z�ky�u��9��~���ݧЌ7�Q�^&"��'�����������O@_�ٵ���Ъy ے��0���{�>J�'�~;�}�v�8ნћb���cP��Fl�NU}L�3��0����Mb�h*����1v��Wj���xp^'֗_A44Q�yE��"b�f���wu[�����x��N����?`r&#$J�3_g��qt�v�����~�w�z�͈CbJ)���`��T�����e��͉L�N7�4N)��-�wք�z:��e�о(x����d�w0��̺@� ��g�����	� L=w�Y�b����O�6���6��|�h{G��BVk�u�,��Z���xG���PM��S�xd��ׁ�t���9�����8QǍ����W"�T���6%�o5�}	l�-A��|�e6��;ВD��j�Ku��C"h5v���0�=|�о����N�����<���q��&�w> �V !���<����B������뚑�_G	TE�Eo�b��~�[�m�!|��E�y5w��W$4��^�f[3=+C��Aے5OЭ��'\=�xN銷���c�r.OO�q��v;X����i�g%F����3�.��\��ӳ��4P�)v�nݾ,�Q��^���_v_��Us��*�l�<�>�m�6/����t�9�y��ϩBD��=�@�"��g6�����`65�������q��iq�@�B"	�Ƞ���vs
��	 C�\��o�~���2 ��r��1����$ZU4��z�L����<�Y &ȡJ!6�JW�����[)c[�`F"��}1�M*�A���뷖 ��Q�V��n�E�{�6�%=�'���ΙiNX���mwë&0SS����Ӵ�1�;/�Cd5s���|�X�� $Uo* �C
^���ӋN���f���e��6��fD��'"ܸ��~��׫�z?;��ð����ώ�$�i��W�=(�[��ժ��g�@�!Ԫ�8�C(�Y�""�ɭ����Y�h�>2 ���BW.�����f0)�^�ft�f;%�q�ɳG15d�>�]�-9�?�f�
 *���5���s%�ڌPk5 f2h�#  AZrڃ��mZJ@ "a�����*RSH�0�4*[�\[��#���c�b�z��9��Ds�-�	�޼*9xO�_��tc�9���³n�N�+-����/ ����R;��	��U0�Ԛnֱ�-�v[kn�=.�<޶Y�}�x�*�6o����/<[j���QL�^��y/�nYBcܫ*Mӎ�S�� j׭iz��|����I�߽��� m�5���� 0`L�Fn�&�4��;�)W�cǳUa�]���V��3'0p$����@�2'� ��*��!����:}�C�õ���L��BDcJ`jZ� �M�. ��%�)���xb�_�ϲ}�th��:Mj �J#�Rh�ݯ���#�*�R��߫����!�3�͌'�M��-g��]c5�)MMLk��*G�O�b����q<"q):9/���#`֧�@�5a�x��� ��؛7~����wi&4Ҷ����P��_������5#�\�j�ї^K����CI�ICC��uݪ�&�nF�N��Z�f]�-��Ww]mav�@~��r�����$6�y�YKwKm06h�S�^j��y@jU&R ��U�M�~������*���#q���X�%�"$ l�N�~R3 �諪�4�frWL�:ϛ�Aӵ��d/�3"��N4��\ֵ����O ,���R���V?8icܸ5�ɲX���h�6|��)�XG�U302RRT#�S5瞨j�{�"R�TD�$f!���Vۖx�!E�P�XT�5,T��B]�O �X��g{\jc6̴�Gv8�|�4��[1E�U���}�~�L���tzv��M��h��8m� ֝�/���b���� ��i'&DD�fS"�lk�Ћ0�)a߶��Ɩ�e�N�P���F��a[�����x�ڪKӹ7P%��e�0L ���V	��q�z��T���$"�[�N�z���~x��A��Z�	�N��!F,U��'>A��J7O ��.�	�~���?01�>zX�21A�"�s�}.`w�IB�*`R�&���:K:M3c����x�������ĝv ����*j�I��l�����nv��p�E��P�:�ǡh���s�kV���:%t��F�c�EGD����u�hh�S��T��l	� �ot;�?؋}S @g��E�Һc�S��K�b���{�l�q[�[l�mS;}�<��1@]C�� t���w�a�>�7i|9!{=N]l�s0���Mt����a�d�$�g0�%�"D��u��۫���Z�Hut��1��Ts����	)�'��} E�u:ߣ��zD�R��j�*`5f�O�1M���S�8�F��	����5��@kk�3Fb�̔s)�@��-�J������ �云i�_#UK-�¡��E*@���+��D���H��X�{���.���v!�H��g�"�hjB)���`pwJA�@L�IOD$��3�I����������jf���QE� �w����C�����V&�=�mje��@��i��UPj!4
��&M��nh]��JtDO��̊40բ� jE��0��x�� -i�;&vX������Y��G� ��]m�#oѾ��ơ ��  blc�Nр'2$�i��FV`�HD���Lv��30c�>Ҧt �O���A�&h!"@ �@���z���%�,00�l9ʞ�:\�^Z���ݴ��RH/�0 ��P	�1���~�È��N��R_�1����8����*��NBF��W.JL��V�8�!PG�Z��1r4�i)�g��\0C��1�Qh��G�.;�s��6;Ԡz2b�bC�>Џ��:/8�Nr���4s@�/J/�	 �����~ .�裏�Z��im0�o��y?����ݖ���O����!����U aa�*RKA�>��E}ٴ���B����j�(�nA�z����#:����6~��#1I��*x�[�a>�ʲVSC�q�Ŕ���-on��T���ڱ�ZED1�v0�oxSC+�9�頲a XJAĐ�j�Y650�;�UG@���[U�"�8����\�"b�`�qPk��)�^*����9�7{<�q�"�l쥏�λ�qT"���c���L� �ZK+C)�a�*����,p�۪���	s�"Z
��ؚR�8|�dt�:|���!��'d�Jj3'��4�
�z� ��SV����Bm��7w���.]*���tEl��)�ck[����jU"��*:�ђ���
�vm-��F�>-:h^�k��"!Q��̪Huo$�ԜNw��%�e>-p`f3 ��-sS;��[W ��1K�l�	�P��BL�H�E����JU昆�
��� �.Y�����E�5rZ��w�PjO�04%��[��	!��!$u+��bٺ�#�-��y���qK/=�Ir�{ݢ�=2]�C�� ��l��*����$��%���y��k%0+Xpuw�3w�B����1�RJO�A��za�d1pz���*����!�ѩh��44f2UHmH���;
�j�������&���Y�nIc "�|_�J|q��,#h' ����*������I�9��R��W��U1 $ �y�u�\#\���[�T�ô�R�` �n_��Fc� 黫AW&^8q��Je?s��E�
��(4.2�����.)�a�l]3 ChI!"���Ȏ�bKSȺI���	��
 Ĕ�a���'�40:�9x�ك���@TG+9 B1������!�V�b���8��8�N��3S���D7�W5A]7b��0��܇K)�>y9���zBB�Z	�8zDE 3A4D���7��1-P�%B���y�E��I�B�1N& R}hM.�C��� �?U}Y�#Ǖ�]""�P����XY�_������A�dEv� 3"��Y���<}�*��{����Ӛ���P�G_��rc �RT�K?>}��� 8���� '�>X}�C��'v��׈��\.��9�b
�ؘ�8;:�FA-�*Rd�3d�|DJG�_��f�L)3 ��)sι��%��qo�O��};Q�m$�O��w0������>�rP�.�)�YX�10��Hͻ��:���|�C`-8�TM��� �ĜԺ��A�S.9��8��zD�ꑧi�n) pk��������; b�T��SΪ"] 1�U@!�D)E�. ��tt5[d΂�Da��a�'�00R&����; ���c�EW<�c��⭋�m��`����!�o�| pW��ڍE�͢�U���*&��@��)G}�!Ұ��0�_4$��P�!�1|�X����B[���L]�wsJ��jǽGa1�` !\`��:�Ԙ&�c%)bD9�/j�Ď"��֏9��	���Ӄ:�.�XF8����F�h
��#4�RJ]����q�9��Tuy+1X���\L<�fИ�᰸2ё�ԕ�Ba�4���8A��(S�H��@Q	�� {"EH�>����u�Mٺ�c�������F��#�m��u�#���CW��).>'s�&)%b��:��#Ct<�g� 0Q%�W5@�Θ��%l'�!:��q�y)vX�h$^)�\�PD������D31sU� �B��%�X���F�"pG϶��9V�86�X5G�[X�� ���an�(39##�~��<�4�(P�1@X��A��>8&)?R� 3y��D�2 ۜ�i���R�袂����<>!$
��#�	A͐0�/!�@�l��*B�A8BWrιd��6����qp����u��� f콫jX^�Eb��>"Ds�.Dj�ُ)��LE�->������ Ĵ�t8)��<O̩�nj!�C�`d]L��RAUM,:��Hn>�
�9�����.�D���	��)��� �qP��;����/��9�ʑM`���
x.��|��R�)Q7ħ��YS�Ήݻt(e��	&ґ8qVq$J�1���)&�J5�|�������Wc��z�=�ߧ������)�d�
�'�.�C��C�Ov��
1����i,=fЛxo�+qk�b�pЦ �3%" $G�N]* ���`&6��Q��E`Z]5U�.�P[%�\2��޹s��[W��KJ��Z�f
�V[\W`j�E�I�iho<ױ��7�P����oC�o���L�܍(�'sd��1
~�t$$�����B���h��Z��9���w���̔0����֛t��s�
 �����2 PU"L���1V&}�]U42,�@U�Q�k�":��옌4p2Pu�!���9��Z[�M0,� �m;8���}���TT�PM���z5K�zo�ۻ^>nՀ�A�ȆP>��F�����;���\���.L��"��'$�L�S�(b|RG�zc� ���|�;���)7�F�.6<.9!�P��z�c��f��4u���9����T��U�8Z»J��7(�?���Ĝ�'�������t ��L��.=�p��qTk8o���I����YŽ����1S��3D>:�7m ����8%&G�FL:�h��0jtpOD	
�����YZMMԣ�$� ]$��wNZJI)`���p�,����pVE5�9x� ti!rK��Yd����c��,�yQI��38�h�0G���4#3bH���;�Z ���8�qe���2֍�'��Sս�1���G�Ll�T��MMK)�<1���:��2���bش����uD�癉km��̦Hfn.Hdj`����)��� *�zd�J���(�Ŝ�ջ�8"�m(L���C��@z�nVrAdQ�t�A�115A�*ڔR1�Nă^�p�ؘ̱�c�c�qf`�������1�D��M���(���Ш�HP�����$;�Hy�`:)�N�b9'&t H)#uq�� ��@j��tt�e� t�Ā �����QU�$"��#�� )g"$�=<$��P���}�E+u�3k�]�12��)!Q�� y�c�B��2$Ir��;y�bZ�����eȈ("��1�jU���!u ��r�I�=�PfJ<��*A��8)ԅ9���2 �#�
�"s���q�<Ǝ`
5�n0>nd3�o7��Rbu�(�(Ls��3 �}|�EH�&�@t�E�ݐ��;������U�Dd�"���Քs���!2!��+#P-88��p�a��=��u��t�5��Sss�͵���c\� b]� �������Q_�Xq�ɴ�n����@z��;��
&�}W7 Ԝr)e���5�M!H;Q�c�����T��u���e� %�VP� ��f*� iTo��(���f.%#��+q"J��\6���		��&�s��ʐU=���!8ֺ�T�8������n�)���n�f����1e�I3)M�H�h�����eFB s�癘����f9��f� �뇭%�P��m!�U��*�\2��v��4CO)S��7���i8�"7%Ιݽ��,�h�L3~"�#U4�B�ED�0�4,������<���Q63K)!�X����Q����S��0Z��B��x��5�Ĳ p�9nƉ	S�KC�C*�Q-��^k�R&�C�Z���C�wH��`d�ś�[ޓ;LS��5�����hJy��:�4"�YM[knΉ���9b�=�	��������|��4�uW�i��UDcn�!F�k�IUU�l|}0@<\G�]�1R��팸c#N8��GCeL��SQE�1eD�(y�b�x�f�oW���AT  `m���J
!Lo��*�w1c©L���!RN9��SN9�i���L��꾇N���yJypk��g�!���̤��	IU�"0�T��3���%5%���YDz������k�����y�"J��xY'|{{}<������r`~%eB7@b��.f�W�8�#�����!��\������G��I4!��CG�� 8���m��q��@�cͣ$���)%NĜ���1qFB6B��Ee���z��H�dFDE[4��D0�`7���J�UUJ)� ��)B+aW!b���r�S��K0�1=��R���R��1Xs$�9 �1� �XUL�S NS)�ܑ�(�f!;��؁T�		����>�*&G.U�������k�RR��f"�h;bظ�����)�t9��"���,�H��Fa�:&]K�
d�ҵv	;V$������V�I!��$*������,�_J�%4��v���QC����Zadd88~.�*�c�mM�"�;J�f:;\Y*;"��P7�wN�E;���]�I���2O���̜���luG&"骖9�r��Gʨ���hG�y��y6�Zw�b�4�JH})��E�4%Ή]]�(�%40�t�]�)"����P�s^��M%�[�K�Dy"3c��	]�H�f#�d���r6SWT;���?���� D{|v0��iP� e�N�	���|>�2�V�ǣ�iYO����v"�)E@���u]�'�Qi艙��>"M�D1�e�a�x���z:%N"֚ �2�"ӭ��6t�X�<<Z8h�Qtk�{o�M�tZVo�M�t^�j�Zf�y2������(�\.Ϲ��w�<2dN9�5�F����V��������庞Nu�a��k���]Ur)�Sm��iv�ު9$fSk���<�)q��/��]}Y�R��*�SꭵVK��ӊ�w3E�Xv���B�|y����k�m*���VE��VJ~:�ko�ǝ�Χ���,��^i��\R�=n�Z��R�xs.G�{?���������[om���˩�~�=�sՈ�I\�u�9���ӥL��q��o�<��T[U�S<�)"�m��E��
�Le�@{�2�̃8#Dq��U��7�*�r�3aN)P
p��;B\�9%NF�"�:ϜRo��8��r{d�X�K�˺.�""�~�Vk;�N���D�����v�%�i&��[ȼ�y>�k��v�譋J�;���}_���ڥ���O"������r:�����\_�}۶��޺\���yݷ�v��SJ1�/�Dv����L���� �Ą�m�Ƕ��T���+���DC=���tr7!fS���ĔR�]T�t:-�J���m�s���ih9��c{�o���u]Uuِ߫��ԥ?����Ã��Zkm5q"��j���	y]VN�xl���<��<�YoMD�8�N�i�7Y�e]����2O�^���Cz�-nL�|~�������S
���jJy��!�Q��B�=*�k��`���Z��r�e=-�����ښ����T����.��˵������E���k��O��׷�������~���~����q�<��/�����e}�������/�2����z�,�ҥ���~|��L�Ut{�S��'Q��s��	 �m{<����+x�x,�r~<�ǖs��BD�@T`�A5D����<OPPΙ�U���Ezo�Pʜ8�*��!��
SN�e�73�S�)ۑc4dF�C0M%�����QE3d�*��.��/m�߿7�2U{l[HmI9��D�,e2�`>CEm�G��1%N��9�2�M��R�P��a�W��{�y��G����H�����ۉHZ�; FC8R��4�R���t
 $�<L]8lF�7%�i*�L��H1��y�����Z"�A(�mb0������=%�:RƉhtI�˶UU	I�1VZ�!{���%��������������Z{k�K
?��]�#T�u%J�ָ�SΑ `�ܥK�u�[��;BZ�UE{��RL�7!�D��tgJ����D�	8�
!�R��������3G�N�z�tu���tZ����ћ�<Me����?���NS�r�CJT#�g��e9�H��XZo�{�9�N�i*u��U3K�81�Z��f�T��������s���~��!h���Χs��"�!$QI�J��2"-k���������6D��������Tk}{WUJ��V������|Ω0��:�ٶo�zz�r�����~s�,�H����?|}���[���o�������L�2�)�\/���������ח�����ۯ�6M����rJ�ƚq>���|����L�r���͡�H�</�|�U������s=�T�e]z�]zɅ����t:]�����㱮���˾o��}��i�E�����rI/_^M�c?���ӹ�m�k�|�����?����p�Ͽ������t�繷�D�t���;���ʾm�,3��n7U�����{W�\.���M���t�)�s�o{km^fsض-�|y���m[�e]����TJ	T��r]����պ�V&��n��m�rN�O5{�}�����|�޷Ƿoߗe�ᇯ�m����z�=4`�K�)�.�v+��֕�⾙�	���f��zrpU�}��6<�(�m]8���5��˯������r:�[o�4���$N��z=d^*��:j�"�p�!����[%��"�)�X�2��2�X�UM���U	�Rܼ��& �rr�Z��_��sʯo����i�k2G,�S�<��<��~^����߾\_����/�<�=1��?�˾凜�����{�km9�/_��[����\��yR�����?0�\���8��t�����~������������4� ������>��Z�q���E��-��D���֔��Q�-ݭ6U�����?z�����	 D:3�ڶm�3��}�/����‽��6"Z�%1��Z3��mj@fzq�]�1�O��t.��փN�V5��	?n�wN�HS��p�۶��Z�e��}�c f�e]�2���.˜8���{�>?_.O�?����䒃�b����,���_��V�!�ɔ�2/�$�[��K�J!f>U=����:�������<��Ժ2=�RP�(�����勹=n��n��a�����������������O��׿������_CN�����~�ˏj�_?��������ۯ�:�<����i]������흐J))�Ty}��r���ה�b8�l��x�����OӜrb� ��D�?�ty���̤G��p�bݷm��]���ׯ�4��C#_�����c�(�ܜ�i�V��O˺���*:�K*�������YD/O�L��&#�?E̗��K.�.-��sV��c۶��K)���|~2�mېp�f��o"��a"��RJ��o��s�yY֔XMUu߶�'�b�}*e=?�����/�Rr�����(���_�e�����o��ٲ�e*C��H���������?���=%O˲ Bmm�vU������z��۽���MՖy.%y��ID����lf���d۾��z�"��DtS�<�O�.3�̦"�̻�q��F��นO�L�k����f�s��^/���ƻѹ��    IEND�B`�PK   �KUM��M, W/ /   images/88f9db7d-1b4f-4095-8375-25787367c0d5.png�{UT_�}�R�@�hq
�	�V�h�-�A���"ť�-��	���C�w'����}����Z3k�k͞�3���Í��R!zJ�  ��*� ��  ���Ǚⴷ�|WUC �����E���WS���La�dC!�z_�$е)��8[����9�J��pN�	���c6�ޓ����Y��Z�X�*f�]9�B�x���c��[�w�PQQ�v����^����-m�a���ǡ����[P�S���k�6K�o�o4�Gϫ�Q�GȬe�������q:IԬ�yL@�c�����0���2������dђ��G�v˽ �D,�zQ��ѕ��!��m7�|�\"ec����x:�D-��}�tT�82���;�2�].mZT��E(m0㢥�M?�}�Ή�ÀYG�W���K
�8x�ָg�B%�ۆ'�[?x�Q��T�Xg����|:����N�)�}�������ϋ�����+�±����3�$��� /	��-��?L������r�ZG1W�#��	��i%���i�mp�H W_=�mH "�:� �&3��Ø9B@��L�Ə�0�����T���o����x|D%��݌�������~�l�A5wC��]�Wk�ȳ�d��#��Sk�ֽ�:g�Kr2� 5���b�_O��c�/������{#H����N31�	���-�y���Y7�/�`w$,ಯ@/��7r���>>7�\���0{���Rϝ;���W�VяX���hk�gs��Gn�����HO!�ùX+���3C�dK�V!X�%�il�^1c��375��s�G����)���_g�l�h�*ʳ��
l�{�&��<4o�����L1�t&uQ$�xSf���?v�Ԉ��c�(Is��~�d�U��l�0 fff�_���ftj^���!�	4�r��U>ʺ"�,IG��)x�b�m`���i��������P�S��~%m[��E�^�N@v�Y�Y�����^���~�	U�./P�_=yN��Us�d�a�7�dY�r�u����(�B����y���f�6����_<���d-)�[5�Q�)x㸚+����i�3�4����a8�H��;v��?���q��l3ث���#�]�(<��>�3T�B�Kla�Xf�{���P��i*����$�|@�j?�HB�N�]��ޜs��&B<��ɢzr�wR�w��(هs���������.��N(:�:��F!�`h}�>�����]g���W0t�a����X|L���o{�ck�roC=(��ų]%r]nI�C��n���]�^��x��H��G&Q/s{�a5id0��i��s��b|��� ��d�Xv�k�	���G[[8r֕p.ܡ9�k���fd*�*��H0B����e�g�	�gr���N����3T�US%W�M�/:(��!'�*s��#�I=���0Wk$�2U��H)
`��%�W{�b#L/p��
0�Mc�n19�ӔC�ʍ��0��#�F�cp2�GO��+q���&h���T}��sTȣ��L-�m��.�nXZ�%���_��k�B��qd-2=uFk�ѿ:�lZ/���20�{��ɝV���9�⃃oƏ�^q����D�k�Cx�(�8X�1�G��~oҧ�u�`�ݺ1)�E�����G��O8Mo�>���}E��;�w�i�%P�A4H�G�T�B��Ł���&��%¡��%)K���f��yÇzx����������Q��&�kBV�T�*���\I��Ckfn~��-��1e��&Ӂ���/Þu���Dº��(�}�<�	���G��W'e�{����/%�'�z�o��m�e%����/W0�.DG{�Z*�z}�6��Z��h	�+� �yU*���t+���"v����(zz�� ����g��2�6z}��]������B����F���G���^��N������c�(���%s�n����������;��d��2 C�������o����ק[�:t���<�D�����έ�V���v�h&��k��>`�j���]ʞ5�0s����԰� ��c�����*�u`,�J�g7�ps�)��8�� �:�<���Y��Ơ�!3�䳝�����=druM�Y�(��,(��1Y�	�#���XuG8���A2NDj��w���7�g�9H�����&UL���t]�
oNOu�D�m��a��IN�6�h����F �J��QICA�?�+�c�o�f�ô._�D����®��N��&�d�.�Ψ�K��Ļ4�+&e>��w��o5Atyi��,i��'�����D�]�1�Թ��PV}��ߚs[i�Yu�o�KtH�H	I~}�'� �>�w��H�`���w�5j�A��r�Í-Q?4��4�6��}<e#J2.�/�����x��T8�u%������ƌ��L	IƤ.^�t|}�m��N�9�����'xv�rt���q����k�����	�����G�m��v3��H�,X`7��A��<t#�x��L�S�fT��`8���~�CoAo�ЗG�g.c��8�q�kz�F�y.��Є�̽OB~�@����2�2�/e��8}/��@��/�w��S���6�=�C��I�~���uy�7����$DM��e@����w�~�7�u���� <.�����iU�Yb�x����ZA���e��4/��?�Ǽӿ{�3��=��FC�1~�MR���Т�c�	���}��J��\Q�H.�1����ې���;�I�
׮����7n.{��|�+�k_��0M
��n�|À2��������Wee�~S<c�J�Ic#�߫���s�~-)�lϝ��;-ڈ?&U+|���U����o�;Ѝ-a�p�
ᴻ6a[�#��JU���)�<�z6��^���E(��TZ�\N�
�YyY%0�$���UM;v�(������T�i�����k��;�:��(��\)Q��
�{�αeTo�@3���mu�����,�ñ.ށ�­$��4|�s�;�'56����G<�v�[U{�@>�E�����(�gH��fc���%��Ns#�7h�w��C�Dw�Yu�\;��>���`P��̛�m>����P��u�v+�Z�q�#�a��nm�t�}���Ƥ�+�}j�����ܿD�'��S����st��m���o���=�`R� �ͣ6{�S����	��N�i>M�~�~�JE������k���k�U�kw[����p����:��8������a���D��ѷ�q��}��@OB�a�v�h�#�Os�E�(r]�0��[��*t.��!
�d��e��E#P����[�]ձ�P���@Rl.x�@t�FL�%�1iE$��F�/FE6|XB觾6�d��$Y2D$���؞��w󍄰Rf����N����X�x����ϣ�܂�l��2���Y������y�����V�.�#��$�Q!����SN�ϥ=ϟ�b��g�kV��]s�ԭ��>�i �%5v+��&����G�G�j�ٌ]`�I�.�[�M	��gT\������CD����UY�~0w�X�p��%K�AtE���1H#�^Ueإ�xN��;�].��H���ދ�Fe����˅pD�n:_3��*��kiH���ϵp���?�F�� ���._;^���� �1Y�d:j6����������o�~X��.g�$ߵ�z���d���]�;�w�E���r����HKC�@:"V��f�x��W2`ddzN�G��׷[����~��R�=���$2=�f�O�͍����/�6�dY#7�,8e1%I��~m����mm�ZXN$چ3|Z�ɭ������nDQ�
�0��K=S?k["գ��!v�G���w9���I֘�g�\٧gN2r��4?{Q/ZW21�
��<;�x�T��1�\i����&��p�ᮩ�pV��]i1�;�4��г3i�m�zB�|����R!�����b���ବ�!'D:)օK���$9�^�c�����87.� [������,���c6����C�g�}W`��IP,�}|z�E���L�����z��G�c�?�!�Q�)b�	�]��ނ���o�=��D�ֶ�%N���޵=�*� _ߛ�u�����M���z4hY0�]{���6�nfvr{��(n��&g��T���W�7&��'qO(1�^�7�I�>)�����q��m��ؑztLK-�{1rn�"�o��0�i��d:Rd�������������X�+�w�����$K��W�g͜I]�y���:[���PZ���k$:�N�[�S��[�q�T�#�� ��#�U��u�h<��?�������ۈ.������l�������ő8���^>��儩K�.V ��p���� l�ʄ��V�|�������@��]$����b��Q�*��Nbp栣I��S��ݒ��j]��O�"��ɃL�Ѡч�����j���`s}[� AQ̝@{��Pê,<���6i���Ŭ������������r,��ΆH���tq�:��\(ft�V��@�|59�vT|��B4�/Q.�/d� @�*�^�~�m9�it��L���Q��(
�f�o tɰ�0	?�_5*���rQ#�Rx퉛� Ύ��b	<ҿ?`���z�N6�r][�x��:��B��]�7����t�)����$��:�p�{@�*��r�o@�СU���Z�a/d;C^yj=q-!ӒY��ʉ�4��o"�4� ?�ǤI�����hs1�K�pvu|9��Bt5c�V��7��
>�j �w�Sr��Y��V@��IddmZg]�#q�E4�#"1x��V`I�%<* /5Nb Fl;כ�wTՕ�#7ɢO~O��G�t����^μ�ʍ��j&ywe��tp7f`�3���v��~`R�nf�N�@�2veM��`�Y�Ǳ�u5~X�TN��,|�A�����4Q�γ�d���s���*�ۓ�������f!eK�eC�,Ɩ��V��?�oV�?,��X�r	��ˏO8Y?KpR��Zf>��g>��}��u����{rq���Jj��BD��.���6�.�y��S���/y���.�3)���?���嗨߈@J#�M����]
v��j8�d�j�8���A��Zo_zQ2I&��>&l,�SZWާ}XdoZ12E�K�K��$,� �M���u5��� \]��1�SO���=H#��0���ؕV�����ʊl����f�E%��׈����K�-�*��+��eִn���Z��	o�����H������+QX5�X��x�|4�hB��xb�ts�������U��s�����#e/�a���5n�\�r���x����>3�QbE������	U������9�����/�`��dÌ��P�d鯓Vˢ�mƾ��N9U�&� ��*b[(�zK���4m,|AS�ƔO:$���R*E�>�e �2)̣҇"ѕ��;˭=��w��)��� �� `��>�za�)b�^׏z��o�6X�Zy�jx"��?�Ur��|��J[M��າ�u��!�x�Hs=On���5�Z|��h���[���$h���B[�`%�'J�<d��WF�ɋ��g�}�~R��nr U���;t@�*�V��:�</� ���b8�p�^�ʂy��Rؑ�~�W�����ݓ��E�=[Af��_JM�_�����e��e���#>d�#/��$�X�G�oכH*�Ű3ID2�Iv�
�����4N=69J]4��J?��>y�k%�O��6)�U���Y�f�)���I:+�ǘ���n��ٸ��	�������Gԅߙ����!��x��;��٪�0�U��?Zs��kCIU������)N���GbZ�Bf�}��$;�d��B�a�����F �=�?��=~��r�h�E����!��ׂ2����6���'?9�ı�-+�G����\�:M|�x�Ir\�1�٘m��<�s�k��HK��	�1������+��m��u������V��S7
��d�C��}t�C�ǎ(��{��K������1��������wz�㽪�I����ѵ�W�ڣ��Hw��	%���ŉ�K�
ĝ��|����axg'���M���շ=��}����q�!�_�X�N�ŗz�;+��Ϭ��D�Y:W��9�z�O�5��w�MQvYKV
[��&))��EG��
J���$�����=�������y��	[%|�9�� ��<�)'e���vs瞥����c���X�� ퟝ�����mq�C�qo.S�,c3I�p��'wW/m��&�>�Ì��VX�7(��&��C�(����L�7�k��[��1�H���^��&ܵ�&̿F��j����)h��n���_w�CFx���2a^d8Ȍ߰�"�e�^{�h�^i�8���TX��l���0�י��2ۚ��	��>�J�z�u�#���Ξ*�ԑoTDff�l[� ��>d��L�b�dp�d��rF�U��P	R�]��6�]�
gp��a7A}4pD��{���z}�e�B<�ĳb�#��m��~{_�U��l5
��;�J28F�{��ڲ��u {���'}Tz ���Uu�6>�U[�5^�A6
h�Oå�B����v�(5�����.>��Y};|α���k0����o���idԗ�<K��[�39W'9~��ƍ.̌�Oq+翍�g���l."?��[O���ݢom�!e�s�ۙ�w����܌�q�n�%.��nU�_��Y�`�֔`cy���}j�K#�Cy����1�r�A������
�V���_Z*�F%#�
�M༪�<|�Ŧ?x���2�	歲�S��ϯ*�.�N-=lv�F(<�_�	�R�����g"�W�[��a��D��b s+�K�� ��j�}tCi�KS�2S�m�7�˒��3�,�7�+� kL-���*�a��!�9k�k#�}��0\p�c�c#u�P�+F�o���a��SO�b LI˩��FQ�ط}�	9�!�}�J�5��>b� �x �m6y���h �b����P��ƃ�
>y�E�H��S�մ�@�1��'��6�����EO�75�Ŭd¨#kTXQ'g�'�I��$/�b�n+Q���$�@��U�AHV��z�����3���~*}�5-�:�([�G��Jx<��^�̴@ga��9�w��2�4L�r�$ҭk��X_�"L�n���_�欞#i�[=*��w�r!�8T'NE,���1��Zb�9��4�va�5��H�h�ժ��U
Kg����O�U0H�h^)d����=(�C�5���O����mcTef X�M���fF}<"P5��9f^�,Ф�ko	��g�����K!�(��
� ./�"G���ŏ���.`'�r��Ⲳy��N��gA��>��qa�e �8�FZ�::V'���O�1"9�ޥ�g�jj5�D��4��FR�d?�U��&��V���-N�8��j��(cg�i$�<+���F��c�+)�jf~U��џ��x�r��y.(��6��a�n��>Mw�$ц��c�aAṝ��b�Ѽt��%�qbDN���u�dI2��E
�81!����._6��N�_̏
�G�mf��1{�5�����z��S�L�rF�"	wV`U�[���;���p��{p-��¸��~��d������R���f��S�~�SNg7
K^!轢�H���#����'��)[ge���sZ�|ҥ��{����(�*Y�O�AI��4�ac�c>�_~+ۂ0U7�W��.>�jQB�c,�&���b[��P%y;F�"�B�<#W���~�㐰�GܠP;�<����8��3�5�6��A�?8�|.��|�+R����N��S�%U;; �C���kO�`��ZI$;m��H�PN\�X�*��{]��3/���̑�´��-��o/�����䷧+i��v�~����L�&C�����"��{+�akj�$~�GGvF��lZu�?o5}�ؘ��D�8��rN�odub�M���o{yJPx�{eN$��L�����!�����%�,�7�ֻ6r��VT���)�W
k�hu������8�ס��q�f�j%�G�ͩ���R��8=x��P�鷹T�]���Mƾ����i�L��B2�Mé���C��ٓH��j�����}]�
2�����7O��)�ޫ���%�y�S�q6�J�2̢���8��yR[��|Ȕ�g�[ U1y���T��B��<��1ӔH���RTȸlO{}�ޚʅ5Ђm�َ8���x���l�<����(�������"�.(�	�ӈ}7��"�D����������[���sJ-����tl����zgnlZ#YP9`�+����?�ĺ�	T�.�^4gY� +� ���/A\
��O���6h�~)9��>�'ߴ̭�4�� _%���V�x�%��Z�_�>[�����#,>���-�D��0wx�w�=��<lrc���30ē"j$=� s@��E('x�NU�G�4�GQ�uhZʩXjs[3�UH��|?�Ǹ|J#0���ڿ��.0؜����c��s��vw1��(3�#&g�P�͒]D `����s�p�n�]���7�n�yU��98�G�:��:Ŷ�����q��
iʾ����M��n��遏�S�q�����@۩�bf��c����l��$�yUN�y���>o^67JR��y�k���ǵ�=��.RU˔�NŜ��S�c���7 2ގ��ҍ�/-�P�M�Xm�E�X�W�_oN/W3v�4%+[Fb�R�+<]ǭ�Qn��"��]$=6���O��Iw4���i����j��`��s��і��)��k`�_Q\��L>�a�×A�_�r$�BxΓo��VҭEg�v����lʢ�,_�erَg�	ʳ�G��/S��%��.o����M�iCg�ɹ��#�H�B��]�q5�3I��OXk� �vh~�כ�=��,o�KI��`9~�O��{3����M��x��{�C����2�Lo^��k�R}��}�k���B8�eh��`l�)BB~�����o���w�7�� V_JdK	��x�hsM$'�Q���^Xj~�B��2�)���gE��;k@@Q��k����L5��J���W)��H��{s�h�n�XkI�`/����»��It�-����MS���&�!���i�[�V[�_*�]�\1��R�ޯ�<��u��$o�I��Q�ƖR�֢Xoǒ���������p`:� �n�����d�=���[�n���?�`A�~oo�_B&�ld�~	W�����uî�R�2�U>]���ډH�i��k�D�wt����bs�wd�S� �O�.�>9�W\�6V�Y�>��.��r��|����>�p��z:�fW^H9�`ur9�y~n<��E��ԟ���T�im�H�%��U����L��	��7��%�E�x��)��� ���K�0ݷ�y/�,�k����ɽ�A��j���+Ο�FL"�(�"���������#}��-�Y���i��qκ�9����5����}W�0F{��	�a���H�P�AoFc���ׯv�a{~}~�z�g/���X��ߒ�"�����`[���R���2���U�7`$6��?�g�Ӓh�	��%Y]���G1���}|���+���\���l�kH��ACK��ak��ZBFG/���ï�T��O�� ?��_*�i$���6+�b�� k���F�km�G��a�j�%�.`�s �p��\fC�>�m��c��E{ѼÈ������?v������V۲���^}:5�g;�_T��0�Q,%�JWS�%�&m<+(.�k�[��TuS�����N�e��E����|� �cdx%�> #�qK�{���~y�/`��!^��N�zn7V
A�$`߷���7�sڇ7�&�c#V�6 �}�%6��.��v���,.�&�_1���lE�A��4�it�)�>q��I��,k���Γ(�����A����"?��� �M�o.nu��Q���v�`�D�O�y:�1��x5�l���\nޤ�Ǉ��6�D&��O�窿��4d�"�ҭ�����bȫ��s�����VkY^�^�Sv<GTj��dT��h��5k�F��19h������U]5��Ұ�)��\�:��k�Ѽ~�NBJ���E�J�/�����|���[j�_θ\߲c��q�>K�ji�9N�L�w�D�zA#ȚN�Z��FgC,�_�@X�_��o㻈��7���Q�O��/Y�I�v��΋�����f�cU[��t�b�������J�M�#{X<gN8���!�k(u8D�B�: 2�R� ��MG��GE�ȗ��9
�1!qa6�q��N��cGa��_���*_�[Q�WMg:
a�o
&�a����|�(Bw�$��>J��[C:��I.�p��v[���N}2޾��x4W�3���}8z4M�UoqB�UBV���
���U���.-���-����˂�G�,���r�_h�����S�ۤ �Id�G�`��i��m�%{��G���g;�w�3�ߥ��n�+^��4�L�W���N�b�fn)
$��E��E��"��j��s-,��Tf��&[���!���|��u޻ɾv�+9W=�%����6����������M��?���U6>��I��4��ۼ�h����AA�G�甠Os�3�����2F�o��{W�K�8fi��q����ue8M�&n��O�T���4j��<����3������Α��M�|/�s�`��X�m+�
=���>v������i�.���[�3o4ژ֌�f��Ų��$[S.�	�L]��n���/������c����z���C�СI��^��� -���Azn����6�%��W�W��&F=��-��TWF<3�y۶E�'��#m@@'����I�a\�W�=*�"=����0Y�K4�i ��=5�K��z0����v��'[�$�4����,�2���Km鋢����є,�礥~-��Zr�\@�g .����G>㥽�K��U+ԏA���~'�V��&Կ9Yk�5��8H�y�5<�Ե�f��F$�m���ȡ����@��������L���sy-cw���r�(t��, 7p��C'F��r�%7F�����D�+�M��_ɓ�H>1�`=P�d�P�a��_�=��4�;nw�Z <��7��{������=�J�_z끗��%`�P�\y'����K�Ϧ�|L��׳b�~n��n�^�$�L�%!�aĵ<���
It�J�`H^�����1��>�u[���nn��Fǃ>L"°3�émJl��
��h?<o����ۢ�,5wlZi\UVԷ�Ł� ��J���2Dm�i���6������Hb\j2'���n#8��+9���U@7��B=�&�F�eU>� �猿I�"�3q}��:0�A�ꄄ�����u^-c]��A�����ړ���`��̹��Pꓸ�߄[>������N��5կ:�'��MN�J�<
���;��.��PO�7���>t,�2�IK��nG^�,hG�y�+X�4�����?v���>@���x���.3d�9���뢨�"Q��se�K��y}R�*Q,�rr3�5���k�yT\Z۲|����y�m@l�f���%��r
�T=���[� �S_v����;�1�^1,c"��R�l{��/�9=Ƣ	���ҝW���o���1�-�8r�Eq�F&�2�
Cm+B��$�G=.�R/Z��F9}۠7��f���!���L3�C��%+��5���bۋ�dˠ��ҁ�_5x�wyqlan*����(�o��+�����]y����Lv���R��?|�J��`7hq}������[�׏e���/a�X�����p�Ӹj��ٜ�r��t��Eqڒ!_��IX���(=�`��.��^}g
��v��ʉ�M��5�!9�B�fZOŊ q�����A�+&�6�����9��Y�Cc�H�����UА!��rX�b���+/�_�^1��C����w��~���6��58q[�R|6�цƛ���$?�|���`�p�g��,���'(��~N��L���櫂��R�e�]�A�.���G�� �ӓ�JZǑ����%T���i�~醟��S�nY�>��M�+�]%V��#E��pԎ��g}_�j�
�m��B(��6�;�a�{�z�Щ�) c�*�/rԞ�ֺ�lF��}�Fg/xʸ?�+Fj�D�k�s|-e_	r0��ް�''�})��O�*��j%��F��T��<�uX�l�T���)�E� u�%�Q:(u���a�&�b����D�v�2���@�jj~r��_�V�V�����N#7K�Q�u?�ִ@���W"{bkyd���A4P,�"k�.bL_��c�:\|�� 2-�D缓W�����hH�~�w�;eS���;
b[�����D�T/�eL�� ��%���5�i�q�˪(2�U�P�s���/��삑�P}j�t6]�����3��w[�-N��$h��61���\�<�^X$����]Q���v�Z©�18�q�ٺL���p��r�.o����d�	�'�׈�(;�e^����lVWr�
8*wy�������\V5���*İ�]Yӎ�2p�Tu����t46ɽkڂ���M&%��X<ζ��A�������#}a¿5�?��.6�\s�X;��v��� `�+�y��`��u�K��V����(��+zD]��e��X�z�s<�!*��Tq)D�ek9Č�dC�z�b�'x��At�-ذh@<Y�O���Id�N��V1\u���Id�����zu����uT͟���m-j�ly[�J��C�����o?�'��#�9uVʈ'0X�	1�(��!Km�Ul�<X�x��Xd��"�25;�ZW�x�_JO$�Jg�-�0�^$��XUpB�e�#�_�`�%y_�~�I)�j6yn��&��5�i�R��T<������xp��8�ۘ����`�Rօcl�.�����KqU�AI4*��s�M5�:��~
�aSI�]��?H<�[wi�� �k�R��:��vX]�ΝlN��׺�^�.X��&��E{#</
Nk����J��?F�]_�9�e�L�J�TV�%q�1 ��=�\�oo�>-Jܷi������ߎa;e���9V�VQ������b<i������)Rh�b����r��b�K���<5AZ��s\����gV
���(9%��[$�P�.��Z���T�G�&Hm�K�F��*0Z��h`�-�,]��2i2�	��<Zh���)�="��_�|�l�5��(������	�H��6�;j��W��EC�03����
%kN7)+ƺ�W��� 4��]�4� �!�]��Ǣ	�\\k���8���zI�еo1�G�$���_$B�-�� R4f�I?�k,�=��*���a7q��8^����$(?�	9���/�Ƕ�8���&.>����A2���V��*W�iZ�F�uNs�;y^;����~�����m�X'�;�f	�Y[ȏ�m������d�6)�&��(2�Ů�`'d��u�C��z�ѳZ������l;�yަ�.7��ܹ���҂1 �����1�fc��1^8����3��c�]"UC Ҳrc-0���� �4�
�F.�ćF��b�1�S��Y�j����pL�����
�$-�����}i��Zl��f]��fm~�f���f��Na��ܶ9s{;K��	��F�c�8i24^-B�_.'\���a1�V_�Y<�ݒ>�Q���^�Jd�r��m�zK�&nFԈ��)�'��¯��B�P�.�+.�gx�V3��sr��4�[6o��,3�����Y�ے��G~H~�l��	U
�I
)��!K:�vqʀ�}aX�-��$���Ԙ���r��������YCZ[���F�P"����O�@_��ec�˖��W�~6q"{��2�ḥ���:�E���ѩ�{FwV��`�������-c�Y8�V�}K�7������5}�~ �1��:�tBY��G�|���Y������������>�~kc�p����dE ӥǳ�lY��r�[��M�ķ9�����N�������{�����l���XI8�2�U;�iˁ������~�m�+%_�M���.3ʳ�~^o]RI�
�h����x�[�b�UQ���n�Wݝ��.j�NDG-ד�A��/s�k���c�b���+˚�L���j�����/��K�:h�S�Wͯ�ƫ<*m�!��Ӷ���3����),��l������g�Mb}��q �_*�(�*�nSK�̯:����gY<�9�$�v�;��ޣj��t���w�/.Ӈ���_�d٥\Nl�?��EE��p��8\�\dyS0�y@��w�e���!V�+&F�M�`W��Qs�L�1₢�Ł:�in�%��ˎ5+��s�isѣ�"�4o��e�t���A$L6u��[���e�R�D/��I�cE�?�Ū����ڴݴ�zV,H���N��qb�o�nx��{��k�N6����f�М�~�v���	r�ށ�QޤN|���~�o�����Wt/�,��[���![���tM�����G�e��e��� ��*�@�?�m��V�����d���YZ��o�/�����Tm8����J��4����oc��4��q<k��`+�	���˝qJ���&��<�갆t#!a'�����_G:�F���&��{Q s�k6��݁�煼�8�/-�N���v��N�!Ӹ�jqݳ"��^��A�ߔv���M#^��V���#��}c�>>��Y�}��Y��?�p���2L13�,DĀ��4�(��>k�*�]���l�󼹸S���YG;G��|�C@Ƭ��%��f��7�rz��n (KLȅGb��	T ����~6f�8*�����m4`F��$3n�ЎP��R��B1i!����Z�xa��Or�P��oUU_^k�w�n�j�jXΟ�� �ZM�}����/�n�d���~�lH�����J�	�Z�lbG����Q qZ��To{��C�}�ݏ���i9�ҞK����
-q#�R���J?�*=kPE��� ���⻶�.!�c"����'���ŵ���'z�3��Iuǂ8G�����'96�`�1�ܰ=��$�?�Z�T����B��ҽ����&wL|MSB�����_�t���x9[��(��B�gq�j:�,C�I�18v5CI?
RF����	�wc�3��cq��$�c�d�O~V=�b ���e��E��(�({d�?y�oH�`|�˾K���B����X�t�x�ǗN��C/>���`�E��\"������۵���� :_~�6�������cU#r��N/��r6ӿ�i�GRV�{\��������������c8�_��f�0���vB�����?T�/�ٽfn/���Ut�T��q,}Yų�3+�)_4������[��:���?�;�e���� y>O�b����)*�X~����r/���8�cU�/G�B���캾��&��$S�U��!�>1Ȏ��G6�"�D��Ǿ]M��Bj+��:��˿�����fʎ|@��3���u�"�q������ڋ3��S� (�~L��-BZz���t�:K�+��oKp��[��.?����c&O�`�R`��
�B�`f$�S;a��U���ߑ�!�����Ug�ԧej��]Y"�C2���}q��3W[�5��Z)�̰��G�υޥ'OX�cN���Z�qܖ�(
�5:\5H�m\D+d��Ňf�J83Q؆��._.G8lq��.,���8�M��>h}�l�W��a-��[T�_�i9F�\�ޞ�h���-�k�L��,�%)P-D(j<(H'B�3�#'�M���*��S��Q�5�~�@�gT5�,?�	��|H�yw^o��rS��
���r�1��@K�Y���hgם����( ��#a�b�壆-�V���XWO2��H�oTK2�9Hp3%����ә�:��f5l������������'�`����*�N.ˎ{�묐vbV���ۿ���.�o�j������t�/@DY�Ǩ�+Kq�^C/�G���8�۸�^�á�iԛ�fB�P�tA��ߎ�  �\�ˑ$s2�Oƶ��ߠO��Z$3�Pu��AxI]��2s�׀��3d��y&Ǵ2�g��|#X9���Z�]�в�Zk�f*��������䝦���6d�/Eg�1F�yFv8y*�O���$.z�c�r6qֽb���K��K������/@пo�n�6)��o��T2��o~~[V����Hﾵ���i��v"C�8v^�>2�O�v�?�V>���ԷK��"3̙� �l,o�d��k���3��}���s�79��&���<a$K���m�Ӽ�d�kgށ�(rp���{���綌�=��_^^2���zz���MB1A�6�0/�������3�<!�f��Ӛiml�]�������1X�Lqp]׵���is0�'��P?
H~'���J�'m��Ժ���'S���"�=�e-9F�Un��#o�~ڨ#"�|n���vN��|>��>��X�Sp�+��l���HmpϮ7�XR�q@��2��[�~��ʈk@rf�״+��B��=P2l����kz,׌T�ց�~߶��{ ���9*����v/:����NG�FL�h6�zS=\��y��{�!x�m^�@�ֱ���Ž�f�}�c#�s�����gm�h�F�ె8j��(��=��H���5�70S<ot-O��Ϗ���IF�	h����v=�ƒ�ɱ$ �]j4�_0�SX�s#>�_V�ݥ�阴� �4�c�������Fv^�0%�x���5gB؛(?�hm&[5S&��>�3�G�j aS�1VWo��^���+�}�ڻ���;ٜ�����	X�pvښm蕷�����=u���!lmd�2<�&�ڍ}���޿e�����A�[\]J̿1c�Dn8`�cZ��y�I$�w�M�'�����Lb�u��33s_[w]����ֳ&1����ՐG=���]��3��a������,2c�̈́�`�gVq�W$�����^��2t4��o�m!��p��d���n�j�嵃��]��7=��g�K�ԟ!,K�6y�հ@�˥�B$UDԍ��n�mkB��+��|�u�y�*���]��Tu&)y_���ϕ��G��KH�4-#���0��5զX�]�d��3m��8�A�o{���r[�M��riJ ��@c2�
Gm�CXmm���m�&I� H�6=�����ޖ"��'�\9�%`�Z!:��J���Z}�����w�I����f7��p_�4�ѯ��r�?��=� 4�i�4U�c�sJ������'����&i>��?���W�ٟ�m���xT�O�`�!6 F[������.�#��T6ǿ��16��m2��4�>Yl-�$Z�T�-k�
M��^�E�;4�1�|��'�my�)��M!z;�-�i6����jF��������7��'�h2�@����䢥9�����.�=|�������(�������%3୭!mh8� �nh�B�Zm����΂ż��15�ϒ�yn��T������OF ����b��Pۄ�k�V,R�<Z���X�5���e9U���E3��������9���۶n$O�	��Q}���s�D �v��}��H�+qW��Z�Zg$Y����{yy��zч�|�%rd]�H3.Y~�!��E�.>�k��&:��ӌ$S�oCQ�
(^��`qkD��l�	��������fQh��=���o��I�w?�|hkF��H�d���i8"<Έ16O�-��(�l&�?Ɓwʪqe��6�B�ioف�DS��:��ŏ�y��<-��Q�/��H��H �в�f̍,��e�qlYJ	V�4OR1z,ҁ{G����P�-�j��ѽ��t��Ѱ���d�䱮)�	��dL�3uC�8��=b��ȭ�sQ�m�n~u�9^NM�P����Bِɍ��a���z���r���	��u�O�6"p�e�Rk���t\kU�[���ͅG����q��걸�x�&q����'�FS�I�VO><���o[�M������|fC��̣𖤎o'ˮ�E�J�|�N�v
;�`�wo\5 �-��p5U�6Ai�[��� ������������D2oՎ�;޾���03�u�jyo�5`�ً�Bq! ��Y{�����l�,�����Pt����(ƀM6��9�yĿ�F�-�Q��g�mK>����`Ub��������Rͮ�K��He=�o�u���k�L�k�w��9��@d0y�N�`>�[�%�@J��?7H�W>��� i��31�ig�]4�.���i��XO��T�j����V��+���˦�{��^y�,��r� �=�7a�*o0I[h] �<�Z#A_ǆ�'%�pH"�.���:�>3�a���a�I�S/o줍)�Q�=�²���!�Ԃ��Fv����v���k��:M���$�L�eiH���2�<]#P���Ɩ�PN��ұ�iU5�{��,;|NO��MO��O:�od4G�^jc��+{OZ�-�qi�X4�8\__��"D�����By^�����O{�}*�}���l�1Xj��ISm$˧m�JcR�LZ�Xg=
��h�'Iӧk��x��d[͖�T�=F�>��7������m��=��U�Vd��zdw�S�읫��S��Z_����#��eԔEc�4r-ƈ�傗��bK5�v��,��G6����1o�P��j֛*�(�ќ��m��9����ݚCLk�b����� r�l��8�V��{�h�5"?�����hb���̟��#��޻$�S�����4��Αm��=�������ߜ]砐���!�tF2���.i:��R����ܯ1˲�,�׵l���Hk�r:�|>cYNXN'��?)1���4�8\�'XՏ�g2�ND�l�Q�����G����F�,�gG��d��Ǒݞ�j� �8h�cD嵽6���m��mC���fy$���:�Q�	T*A�� �6�h���o^r�1f����$�`;ƑglSn�\bN tFf�6��K���&U��z�������:���|�3Ӵ?���������Zn���O��7'kjw�.�)��/��jC�n��c㝷�?�[cX��c�~���'{w�am0?����! �ZṪtB��U�~���!��P����F�]�HH] w��w�� j R^K��Q�G�-�W��{ �Q�������6)�=j{!@Z𠁸�iy�wu�T�ѱz��1�,;��$[�[M#�i ա�3r ����g����������v����s#�rP��lI?\�1�7v��J �k~������{�/R�M�jui��u��!����zO4 {����ytʺf��µi��]�|*u9�'��XքT?VtX�R���}���v�9��9�x��V�:�vhGD븒�u첈1�Y�z%{;귔��_��Ŭؔ帯I��y&P���eђ�s �d��=R-x8?9�`����`�-�3��y����z���k39R��֮����E�^.��r��0F`̕�̣�I?'�1¯+b6�x��l!O��9ps��pK���[��֗��-oX����Wϴ���8���r���b��^�_�{&�8��K�˼��&[��k����r&���Y>Ի�W��wjX\��|�!��Z�"FS���C�c0�!��c	�K'Ć�w�`�� 8�ha��!�mi�I�0K؃�tP�v���e'�c<�z��L* c���k �m���e�Z]��v�|ש]c����য়����v�GU>�&�;W��7��ݓ��l'qp���������i�"Cu�9�)%@:�u��Y��~'��8�0�
�melАc.�a�?��c�#M���!�h�¯�!�8#�mW��=0�1���jV:� (�l�M�t��?�1m�Qk��=��1���#M	�~���=?9�c��2o�ަ�G
�GӤʹ][[j|O���i�RY5����W�o��J��d��#��f�=l� ]�4�d�ҞK:�=N��5���p��0�oc-,<�h�v&㖴�3��0�N'��"2�S~zկ1y��p���e9��|bhAd���zȵ�W�&.�W/u>�F�=;]�#�&4��{�gE��뻲!3 p֞���X�y\�:���p9c��@,y��* H��M��PX��;���y��r$��ŽlERE߄��ر���sR���Ա۪�R��E+�����v-��p��C�81��8�ۤ��ݖYK�*�!-����ޗ6�H2���!�&0��,�aY�u`qX�dTEfj�Z~��a4�!�Qה�d,lH��I��m�wBZ��c���F/�x�U�Z���6��m^�&�orB��Cr��}�V��[�Ǫ�76��p��Ѷ��H�@��Z����b�i@�N�]�����GI�޷��@��6�M�0e��Ce�9����z�}�8u��|{L��nYO���s��L&��{�,�	�$E&���e����2���͹Ʉ�m��#)�͎w�ʈ��l�a��o��	!���P��#���2i�]�Te�̂M)=z����Q�.�4����^��:��]��4�[5J
�&�Wz�����H��ɞcJ�ɺ���+�y��.9��d��qF��I!�#[��}h��fS��V��%��������\
~���(��{�ɑ��,cV]>k�ӫ�_C�G[���n���~o�=�]e)y=��І�n*x
�Ԧ5�g]�~M��X�>ѐ�ur4֞���|�M��`qly��y��,�Xv� ��c��IgRl�ȘJ���K������y�:^�&�!3/_d���I�C�fD���{����w�\�rˀk!�e\G�^�(��n��޴O��i�9���[룚-�^��vf���d�y���}� ������1� �g8��f���A9W�/�lk�)ޯvo�;� �� ��:jƷd��ޫ��y��֔����ؾ�޹G�^���j�̰a��9?�47*WFh��Kp��e:��:���y%�-��k���mN�����}l����^�Ʉ�Fs���|�1�B��?+�,���6�y�-[��S�#���h���es�I����*�!�b"��# ؑ�6��hB"�Lk�L�<�L1�)k���6 �R��"�8e������M��=��6`��s�������#�q��g�����gy�6o�׵}���$ze%�M�Z����׸I`9���ȫ6<o�)e?-²`��'��L�z]SXb)me�; �v��<ĳ9�MX�GN�}�}��Q�s�b J�'r�#������ �D8\����ENe�,<-�齢�e�$�c1��C�c��Mv��v�I��\X﴿����!m(G�<3˘��g�4!�\M�L6���6�uCO����A��S$�1ͣ皊Gh���mװY�~�Yl��l2�89�$G�j����j{I�Cu����H�AhY\	����z-s쌍�l����v�Y���l2=V�/qc��;� ���v�m<��z��#5ő�:bh:֬cO�=o�8�<j����(�QIag���n�+�D��d�F�]t��G!{z�A�-!�$���\%;Ti�.9BS�bv���/�+Xx��6Ɣ|� �ʘ�9�hc���!�'�B�=S�#6�%<D�V�_�	m4l��XTǱn��x*�ќҶ���قO�Kwa be���^*�D9&�'|WM�ҁ����>n�G��6;cp]W\����2e[�v~<eS=s���l>c���i �,�6"y,�"��`B�p˂�:"��2�O����Kx��///��`�`���&�E(ړ�tlD���s�g�ͅ[ N���v�|!  �36�{U����̎W��ɷ�MkV���'%�4I�k����v��ڄ0#�}����Nx*g%��e�{_��R�n�F�9��Zo5Jo&�΄�˽���*��r6�u�؄*j����^R9�r�'�#��	П���=�#�����
�����67��a�fg��ͧ�H��`���U���'#���>4im�4���5�`�~x`p*�p"�������js��&*iȶLieD�z[[��k�]��٬�5)��W���+�s�ŗ����7����{:w�yɳ����a]_��u}�z}���#ޕu]�s[&yyk� �L�!�6�hal�=�o0�&��N n�qk��G�v2xLz�=0z����$�-�Ŵ�,��ބ�!jBV�h�y	~	��r���[�l�l���<�����j�,���<w#��`s��bnyk������ѭ�nk��;|s����R��ѭ㌀��E! j�[60�}�:�ك���^�:ΥǬJ ��`
�^U�6ϘoͮW߿GX=��r:�_*�cLT3}��@`'3�]1F8��X�\�h��|�S'��~��cLٝ3,5P�iC�~D{5@���������1MhU�G��F�i��N}�����o�E|+������3b��;GlL~��������B��z3����u̹G����-؟)�'҆M%��n#P��X��<�� ����I�v����Ȩ@;��l_����(oT�/Z$��H���bon-x�\�9����s屽����e[�ڤR4k�f�z�6>&��	>�����8�W2��~ݹ�}�S�.8�(F3mhw�(}h��܍m08������9G�&?o��W��K?%�&�zK0�^薑��r�Qd//i��s��/�;�>hJ��^�@k/�A$�06%u !s^�#�Q{e[i|=ҁJm���л_j�Y��lH��ȳ�6M�(�����u�lBVμ����̪ރ��z�<N��[�����������9e�ٚI��m����^�d�S$ ��we/����5|>��	� /�E6�}�I�,���͜16S�)7yO�қ���)�y��Oռ�~��:p�뭷�Ү%`���1|�<^F���T����֏jS�)jGݵe"�l0�����MvN`��Z�/_Ω�� *��vg_���qh8�=G��L�l��7���:@V����¡ ��l�f��=��hN��m���\����^��6��9PSm��0�6���k�?Z�Mt��S�s,�6��d��r;�v��e��cm�1ư�V}S�f�c\#'��'�ڦ`��|���������~�������=������~������4�K��%1D�����d2"�"9�?��BS��\І�ܤ��|]����hG7[�fH�S�|�q�G�����&����շ �4�$D�Z�,�w鞺���e蓏���T��"q�������b�V��S�l���{A�fsI���_b���6���Q� 
o��v��[H�U����2���{�M�\#�fJ�G�c�0>G�j� ���=�7�l�'�Uu�_WX�(>�H�yX6kx֬�C"��|��� `Y� �\���ǙR����ՋT+_������?o��I4֝�ܹ�rgګ�(G��3���p���P��ܽwS&�N��t�Ǥ�$pH��Bjp`�D�K�&��:V�eϦO���(�0�4n+�m.5�H�:�����F�|����#�H��`���K(��Hs��K°u�w��%��Oeyd>�����<��$U�kX2A�}��T�����������*)e��J�x�3��� ��aB��t� 壄�Sw�o2qM�[,�Ӱ���d2ۇ��
�m2��-6�{�U���	^k_O� �{d�Rf@�[��3��@�6�/�^�q�va����b�=�;��t�#�wLup��ɕr��f�>ĸj��"7��¯�v�E���`@�P��G!�T��`��{�� ���GţN���{�MlS��ܰz��d��o&��k�mwc�uy^q>��6��t�w����w�G���۞�&�T]��Xw�X�\.�!�:�����K/H!��}[Z�D�y�)�g�b2mQ-[�;!Fx۪U���*�b�Y˪�Rd�h��Hy��*d`�`̂`,֐'{[���`1�Y��,j�suG�m���\4[J�>f���-�=�n����*�ׯ�FǤ�D���:�(̄+����Ucκ^��B�L۶��Sͧ�L.d���ٰ��k^H�=#߱�K�d#�l[��H���
H�gQ{�emO��?O<�7=����G���b^�2:����g�R*�x�cj7�+�Qԯ���>O���x7v�bl6l�⑭�'U���G�o�ߏ<����+[�K^�g7y��G`��'m�e=�Z2����ݪ�Gk�,���(NtL�а,�e��B�*�l׳�EX�`�A�A:�
������hY���'�`���e �57��ReHG� ��5�X��46�G�Td��$�H�~�@2�G�}+5�4ľ�<�1�L= :~g�g�Be�հ�w�_oE240w��Do��E�y�ʘ��u��CR��71M@zS��d�9�X#�N����|+yː=�����rҢG�F&{R��ވ���g����i#��:*g֭`����G��\��o�&/��)9�,�.�����LC���*=B>�$I�v�~A��QR5v��-;�f�|�AG�3���'�T%̶q�~����Y�Kn��ܲ����$�Z���
@�2�
g�F2bɤ�v�q�	`�ɞ2�Q��c�)���{&3��r�8ii/If��\�][�&o���T������Ym�ٕ��?��o9��yJ�$=`���WcDgא��$���ayT���i��Aj���(c�fw3&6m/�8�Iþ����T 3L��
�Ξ;�RR�s{�����
�xgN�9��L��e��{�jh�t�m0�cR�-��2��m��v|��ʎܺ�����p)�^�?76�XS2� ����]^�U�n�z ��Z�
���I�<�Ss��ә�8J#9i���q��o=3`�@&U�����iy�h�1EyO��YV@~��Q�5��wT�T����M��(%�9�C��OmW���u��z]�������1{fB{��~o!�
d�p�gc�'m�52�6���@�1F�sL��S'M����� Ub��Y@�����b�({ߞs���4�ə�d�S�]���}[/li�׫o�{�PL�o����"��+�������e����5pfi��6��I%�h	4�{4V_X��I����Yr��A!I4;)~�py����6�
gBe���6+׫�J̈Tq����}��l�����LH$�q�ห=�f��o��Xg��ppr��y��C�&�� ��Q��z�8���:�g�?��}?�>j�1ιS���o�zx]�:8ka�g\�q]��u�<|`�6��5�#I�/oo��{>;�>)�<*3���Lv\	*��J��t�u���ܴ-�"=�S֋3v�JVSW������s�����vW>
��h��h�IO���i�H��R]Έ.�X���#ة�6\z~v_��s_�@���GE:6,��3ٔZkabD4���
���ꛞی��̦m���l��&ZP���0�Y����#B�	�;���&\o)�@�G����\Fc���{,,g=����u�>��5P���?"��Zݟ]>�<� tD��]�-q�����?ٚY81IR�A�5��'��r��Q�#�O�˟��ί@�ۈ���p�h����F2�u9+P�ϊ-�s<Dy���d�m�ʗ��#R�I���UגU�� �A+g�c��'�#���ה9�	�v�R�D�ņ�ְV3qI�����ϩ��z������T�=/�b�@�ڢ��w�;�]oђ͔��������X-(�Z���nz��ܺ��s֦��91��C�fջG��b�i"���ɂ�^lH>�|B�	`�"�^�tb3�)���Bx��3:�\#����� W��ZOU3nU5~e�\�{�K���'�ɉ�0���BqdQ����e(�����*7LV��N}3�YS�ӧڎ.b2�潢�_l��6��Q�$k��y%��Gh	���C��,ͭ��ҧ���3q��6��;�u=0"���v� ��(�t�,c�0�e'�����Bi���3epͽ�ba2�s~yy����f-�r\hn�9���<ٌJ�����gd6?d��`��s�1�c?��pBTY�"�_��p�̰�+4�� �n���W��j��t��4�~ق8���m��vQ���u�,s�2��EҖ����f�8@��HZ=ɰi�_Ԥ�0Pl�\�ա2+�f��m�>O�7�6 G�E�9��^Gm��Yv�0��}m�wBٜ2m�΍6���֍/�����ӄ�Эm�mm4b�S�M4��dȻ qr��Q8z�vxk�7�C�������:M��M�M�o�(��̧�H�4%{����ҌQ9�L؏k��\n{��C��C��g�͞��Gik�궛k5���gR�bH�ሀ�׈ c���]`�	1~�_-�>}���o01"��<���G"�I�U�����3M��+S������e~
&��"�&s����*���`�R�N����b� Z���)�|�����N�6�R1������tV�9j[*�vU��Rࢅ�h~�`	f��ƤN�iQ٪�ʌW��1-*4Vgk�7�i��o��HN�D�N^'�H3b� {DnyܾS{F����h��ˑNP<�!�b��Hu��MZ�@�Q��[��н���M�Ge�������WϽäfd�<��S�BXG���VgY��H�#�vlTN�amC�ԚIeT2�>G%���ݦ�9lr�k� 2�t����&�l2�.!x,5���x�������ne6G҄qpn��=���	����95y���&�I���C���VR2�t,i�)U�ء�X��Ɣ��3&;��������y������ e�i�c�jشL�[��g�=�ٔ7X��F��zﵓ��0O!��N%4Ԗ	$���э�,���f��D��*��LhϜE�[ڄ��m�>����ܛ���j�̓�_� T���ϳ\[ئݜpN�
������º,0�]���uů�:��Ոﴑ��m��[�1)�d��`2�[B����-�jT�Ơ2���c1$�A�ml2�ʣ�fic'�e��S�SY�ַ���9#C��;�!G�H?��afB�u.ٶH2�vI���l�@�����5t���x�`��ᦚ6^g�{NHr3��i��e����A�g���D�a�cS!�˪K�=�#u�=�`���@�͟ǣ���f���kC��G��;��3	O��3��p����ܠ��s����	�_q>�p>���^��G�#�k����d�FH>ȴ��Ԋi�b=�I1��C�n��D�Fc�ܒ�+9M�,��j��az�k:��k���-���kߥ�-�65Ǎ�I�NY>}����^��}������M�bW��"=ЫOֽ9Ĝt�5�1۱S�ulԧ��ԶǦ�^�# �Q�d?���8T�|+��Cr�(�09j��wFU(�֎�ד�����^�ߋBлF櫖��@�R���e��"��`Y<fP�dO�>�f[M � n4��5��h2�u攞iH��${6҉��PF�Q=��e�����೦�_.W\/\.W\�`���5@�|8���c��-�-X�+�Ӂ6N&��ԗ�!1�^+�zZN�}~�|:��Bʹ��պ� /;��T�B��b��E��Y5��l���N�`̾j摴{R+S�mu��@�b���|��m����:i$��Y�� �E�M�K�ʃ�����̪G�[,LRP�؂� �Y��B��o[��� ���c:��X�^9���OJ��I��!S��
W�7��&�O�$Z�K)�q����=B��( o3'�Z?���,mPj����sO���V�Q���񚥯_~�~�X��_��x�m�bl�
=R�>�����	K�x�]� }@�" �Yk���cH��>XXB��'a�{���T�sߺ��xj���Պ6�I��H����=u{��d/�K��?jWV&�\֑��9����W/��ə�o�����6�:{u/ڻw�5�������*�>[�m�!�#��/�>G���*��<���ޟ��٢jᒨ�������D&�^/�����f쀳0��6���o4�A��^�s& ����4ט��K]�ky��_�c&��H)���Z3�9�E��N��dLf�[�c���ʙ����/����:��B
�z:�4�#�Z�N�)li{ͱ��G$-R�8���0��<�H�@v`�N>�F;J>����{WU�@H�j`����$�-�#{��SJO%0VI�����R��c�6�0[�B�۽�b�����=
h���v?�H��\�5��m���Y�����fTߞ��>����_��PI��F2�W2,p[��a�9�=BF�d�g�9ڷe����6�q�E�X�G@�I�<��᣶�n�P�� ���bm<�F��>J��q ӄ��8Ę��|F��0 BH/,�n X��a���;�1 ��`�[���D�0���Dx��g��� ��ǈ�|��آ#�1�p�948�y��o����k6��F������#{|���l��m�d���y�ܿ����u�x�k���e)23��Q��NSU�����º��"�=X�m������&1n�Y�_�;��,e+�/ga�5�M.:r�SY�v�y�85��Ƭ������JGr�� �o���`N���ڎ�c�]���u����&��Qp���8��������p���b�V�Q��MLЮ�M'���?z��9ϛ��/���O#�yɮ�H!�7��7�je�8�C�<��'�Qmb�8y��1.�1����& � �5�mc+���c��6$���
,�f�rF�L!J>�>	�i#��b��<g��I��6��o��W�t> � ��ҥc��жS�`��f�7S�^��rcx�?k4/�X�I���H����6T�f�H��umO�}��{�m\c���[_�}���7sO8?+4�~��&Ͷ�XU5����ʽ� ����VP@�ԝ�Q�an.Ҕ�q�!���PH�^Ķ{B)i���U�9�=Zn�S��F�_ p�\��2M�6rD��q').���ԭ��m,�'o���j�)Yz��H�1���֟���#Dn�?�|
��%u�4Ҥ�����d	UV`�<�1�T^����gm�V�5���s8��
 ��[F�@�5���@�,"I;�n4M{w�����oUÏ&Kb�6L���H-g���\4�X�hM7d<L�X�@�j��X�LZqN��P�c��?�,b3�����8	�q߸�E����6��%>G�
R�-,����9��k�H��jd ����3��-�����/�>�?�G��l?c���$���*��3ƨIJ��Q�͹v˵4�E��$z�XkJ��{l�)��0=Z>ȼUz�L���YSG�ߒ�STM#�����7=�Ld��m$G���&l�k�[��5�����L�<f�2*�N�T^���B��K�1�ɩQw�A�ptl�4��G�hGa���������-��D��:��@�Ǎ�)+-����)7�� ݷ�����޹eL�zϦ���m�%nrA�{�_e�n�L� ��˩
;Fo�z7�!6a��Ag�߰���r׳K@rUo1+���|�8���ӌ#�~/�ښ�ɶ_i�}�o�Y��ί����dv��8��i�2)�*�x�"�=����,�\��&���|�i2�����TpaLr�	 �g��2f&��4�-��a�u�-z���iwF]~H-8���f�|h������8��e��3�z~�ʆ4��<��X=����;@Uއv>�;rh^��: t�Xc W����� ���`�4�Db��Z�~��@�-X2��:+{�>����!�z�{�eя�0��$��j�\�����7��j��b�C��s߁d���tm�u��J��GG��!�=oLO��s�5?��(6�d���Aה�Uݵ���Wy���y_��8W��s�}?2�O�maL:�1��_���|2�io��r���@��8�z����c���emk723	��46h$�0��Q�i��g�u[u�ڦ�;<˙#�[	�?�:�����Y�f1'1Ƥn.�C� �2ysЕT����(+*�G�/`����H`��k��+-���.P��f�q����2R9(�c�5S��K֘����Ԗm�X~	������8a�K�͒����E&yty3Z�9y�8�4Mj˘Hؒ#ym`��J$��$Vnb��we3ﲓ�������OQ>��	0f;!�p��A��J1��Ui��m�2�Aٓ�J{���d��#mR��s������3��#���*jf�A@3D3�P��i&6ngh�M�z{���މL���h&&��ϖ?{҆Us9*�a����(�4������cu4����j�HPO����6�XB�4��nk>Nf�N�}v�&#Pm��n��bt��X�I��	��5�q*�];d�D�KoRF Yޞ�OjGkJf�Q5J{⃇��1F��}�|�Z�ɇ��M�?��Mz���9XH����c�MG���{_�jP~����#w9��#	�h��Jejm�Ʀ'�XL���j�G�ى�f�w}}-�����n[�G�@7�C��k)���	���kX���G �'z �]���j��������j���vc *�>���1"��aO�I�_~���#e�~TS5��6����{�[��5֘<��� �c��'G�wc/�y�3��D@�C�@�j�>/	:� �*tnIʣ�䚢FO!�[q.�橽����G����m�j�#I8fNB�1"�Ǭ�Y����Lc��3�����,�^=N�\__�Y��v "MWKL�H�a<b40��|>cY��!�|�@ލ�)���Gi �6�P�)�M���.��#`��b���	��zf���B���	 ��sw`	]���,��b�٨��x�FY�4�����9ߘd7�S�j��HP"��\$y_���N��>�M�v�Y�c�b������r<j�at�2��r�~�|�;�!�z�"��b���$�8���+�6`��LY���1Vs��M�@%�#�er�|����Gv��F����j�\ړv7���1=3շ��q25���+����<����o�!��L��o6D-��k�ڶ�j~�6/�����CA>�r���ۍ_�\��[`]Z�C�R����O˩$w!G�N�=UL�8kJ[?��&2��B,/�|&�5@y�1VG�0�K���X�Z�m�����Na�����q/#t�T2}�n��t���ӽ���h�a.��{;�:=;����oCaQ�V6�����ƎJ��.L"��Q�$��h�S��m0o�q��ݍ����Tm���k�w$��ؚJ�:�m� GyG��N�mӵa7p��vwڢm��]P�LɆj�ll�㞰-�����}P�6R;��(��Zm���on��`7���;RЍ��7��`p~��k��e�m��5H�����: ���q��^�����`]J�n�87�9�R_������G�C@��M�ζ�0��^yκ�<����h9P�r��T���X�]��{�S��~;RG �.
�����.#��m���B)H��n�����6ܑh���1ҽI@����hLl��U;�^|Y�w\[I�v��>#��j:���������Jg۸�d��F��T�ܑ�׾�q�7B��ړ��Ex������R-���=�����=#�1)ĸy|<P��=9����"^��0W��&��r��wl�_�3��4l4��t��y�>��76����{��P�����ӾG˽1�-�B]�y��+�XҾ`�.����Aٽrr
�~���^���W��Ò՘G�O�2�u���,�ZE%+�{��v��c>��4˒���K�f��Rz �6���T���e��!�d�]�C�ȳ��L���,��<�"�����%��w)�FMKv����X\�l���#��2�{Ӟ���wY���׾�	L�n�y�g��q�	�{~�L �S��>���A�g�������GH��=�͆�B'����FX�;���� ��f�R/쨮��r�6_��sj|M*#�+靓��	��.���9 '=�<�����so����m��T�}������,8-V���-�-�[��2Nd��� s���omNlD�gj@�S��4�����6��sY\��[u\:ױ� #�(��c�V�r�F�;Ɣ�5�{��h���p�xX���ƶJ==�{U�o�gp5� W�&��͈���λ��k�Gӎ	���Z.p�L}��=�^��yԆ����}�{Lo'W&��S���b��n�3�N.H�������1ƍi�'��Qٵ_��j��!S���ߔ�c���6�T�=���C�m=�^��j�ĳ���k>J8+�,��t���lv:�I�)��^�$�͐fP1�͆U��oΧ3^__��`-� A@������	H�u>��|�9�)��Q(�S�)�z��z���K�ӹlc�?�1b#��Q��柵فآ�����}f�Lf�	)�g��-�[��s��FĴ�X|�}5���!#��=v��}+��o�� ���_σ7�2q�k��Ź�ci��m�����v�7Oo����ɳ���{����Ɖm���=FMK�7+�u�X�3"Y�['J��ypt~lt�<Z?-���=R-5��r�m��FW�NsV���jq�Zm��m�6�A�3�&ᚒ�y̦�F�9g�h����K��#"=�y�&.�9I-1^��[�:��r��%'����k�nN��-�S~?�9��J��e��b]ה)p]?u�������rΖ�l�����Mj�QV�m-k��FN1���*lR*[�ɼ�Єe-�dp}�f���م���p[F�K3qHVN��w���퉴ݜQY�U�p�g��Z�np4��K�JV�,sc}���-!n��h�<b���.�YlG���Ʋ��{�=d���P:3^�G��kBCsi���@b��4Q�����r��8b#[�1*@S�_��Gn���Zb<��sY#=�Nnә����؉����3�r��6{n��c՜<�e[Gm��G�f��O�d��쥛��z�k2�l$���.�69������VM�Io@=jALm��&�>_>1957�aݷ��W;1�v�i���=u�2��8(^���3;�5�oiS�s��1\1ޖQGۀ� y���[1o=�c~����;f�=E�<������%;l�y�?K��� ��Ƹ�9�w)m4�i�-�-P�yfh}@޳��&���o�pC�ٓ])y���i�WͻB��2#Gc0������1�`{G޷B�9la�˲`Y���_�i\<�U?O��F�� f�1֧�Rv�9���o�v0��/-�b�&O�h��LH��X3�hc���Y�Jc"\'�~�d�
8��.nYp�^aMS`l$z=uS�J�'��A���@T&�N�dn�bRl.��R]#v�X�L��L�=����x;��L|Ic��ȶ��}��%��@_иmdo����Yl�a'�Z����&V;�[ԾR]��qo�ձ�2��G`��|�͑�ǽ{�Yd�(m7m������K9C϶��޻���m���y�e�T���4����W���gSVh�HO��m�DH�[`��Z�s)Z�xyMo3����޷D�^F2��Y���������dm3#�L���/_���?F����r���j݁l�m"[B��ڈd���V�f�KR�{��,w$����}�|8�I䐉( qsN��\�h	>�[��5M*�k`c��n3����ߣc����	<S��b	Nl�+vM��A��Ԗv�-A%?oxO��]�J��GR��'e��� i��'��C��:l��fB���1IM�;�oZ҂�?J�m��^�#��?�e@!�,V��c���Ws��,V�G>3c�ݟL�*A��6Ɇ��k�[�����v?�y�{�K9����^�2bp5g��|'��c$������GdϼlOx�d
���ۯ�:2}��cM�#kjn"��ow�q�S��.��I�����>o��k���YJ��xnqe��W;=��,m�L�=����-B�y��@�̓���{vhr帴���������芊���[��θλ�dcSE�w �A� ��􁲠2p�2����EH����U_�}<�E`��1�l���`�c�2ӽr���gĠh �5�{�����Oq�Q��lB5���쵯w��|�tOhޟIk�CQy$u�gO���wo���1�@��h�<F 3�󇢡�	\^/��([��Dga��ܷ��3�}�H�p&sF��ogRܓ�r�uu�5&�b������R���G���0�r�:i��Lz�*"�& 8�ﰫ�a"���/bl��Ȁ�Z!	���;n�٫k$�� �m���@��)�4�6ZA��~�-4����~����-U	 ��-އM|>����4�g���X�4�p�(�y[+��R�nG��|�҆S�d
�ſ���k�=���܃E�tryT4.���ٯ�c����	��2�����1��m[4{ԟ�u���-�kyOG���|�i(lQU�gx�۹����S'�6�֞��1�p�Z���������O�|�_�|�5G�~}�n���e:��`�̑��u>���W5͚�a���y$ʼ��y��-����T\�=��w� �2�DSߙ�.eDJ���^Po����;ێ�m�b�9л���Y����W9>���e��:��&�^o�|a{+�15ڦA�C��#յ���奰=R�x������T��j@Mn�(m���7��u���y;��D�?jK�v�)͗_�| \�u�����qj��B/��ͳw��|TZ���ך��~�i$p�����AԖ[���������,dFV֡ܟغ��v%�`(���������{��&�d���aYG �������`�n�[��{���+�r�w:���'ӏI��l���4�D����D.^`�����$��uFx����(������z^�=5�5)+�g3>�wl~6��T�	�&��N�1��뗣0��6F$ggM���&\�Ѳ�)N�Qk��e{H[Q=������9��!�1i"
s�=M�[�p�h}���8����O�;�~�*>_c���+��{���
�W��#� d����{B3���i�dV�Ҳ�/)9FX��h��	��}]��5.g	ڲ��.�V�S���p#�c�iK��r�Bd�g�X��[�3z�T�G,L�t�#'OΈD��R�q��ߏ �{�H��Ɣ�wB���v��� j�����Te�����5cL���|Σ����zw3ƨ�27&٬�3��(;W�EU�3��U�s�u�QQ��Q��̙z�*�[��z�۬�K�.� � f��o��(wS�MJ���s��[��̱�TZ{��R���9�@���ȩ���!�y9�uGX��9p-��)��n�������BfX�U���&��&t��W�����Ne�=�g��̻��!�5zޏpj�6^.;��Z�vR�9e1�5R��'R�yҾ��ؠ�ַ����=��b*������5��d�K���@�W���qTE���Ek�6�3�&��Wm����GZ�H�]J���H�!�����������ڔ���+�������r��i�s��)m2���c��dx�hZ���b�d�
�V�)gY���ܟ�����c�i�4_^^`�~]S�jG������p:-8}y���3�G�?6�:��ޱ��27y��o�@�Ηu6�Q��F�[0f�NR|��ca�v���{�>�ʐ��(H���xc�ޫ��790����"�D+~��⺮�t�Hz�R� :�l����Z����)^fr�����zC���z�7�|i@�Ǩ�vh�� �G1���1ڴ�~;��7v���D6���60����#��Χ���9qm�NV#Yt���~�@�ۤ��%,�s��H
��L]�������H�� 9���<bae?�������J,e���a�_��o�s"LQ���1!����7�����h,��x}�"�d3��A���-��	���Dx�Ϯa�4 sVzua��<� X$��&b�)fi�݅Gbr���L�v��k��Ƕ��q�]@�_�?~tbz;"��m׊׽M��hW9�V���M�l�����&Q���b�es,��f���v<��cBn��}s78z��J����uG��fFv줚�o��֎�6RF�"w����մ�����X�z�S���D.�4�e٘��r<:�m����2�8��g���O� �"�-V���0Dd�ޛ�m����-�gЏ�`85��|+�o�� ���y5c��V.Y��5i!��)j?�M���vsN<���=�5���(Ez��J�������g��5<�ӔK����YP8�H!+z޵�Y��C7�Xpd��s�d{h����V�c����F�D�gcL�v�n���KɥU{��k6S�����Ql&�Au�iWa{�EnX$�8z����}����xbk�#���`�"i��*[��es�В֒��Έ���B=(���y�M",6`��vHs��K��6�����vN3&"F���0]`���7{-qWa���=�A�gg.�|j�yD��1��O�\�y�����f{}О��֞@����TX���qne0%*���٭���b5b�hᡸ�!�Ƨ�r���Y�x�>	���j���Bc8�6��ǔn�M�V6��}��5jG/��{��{��[eｏ ׭�벿�l���%�N�y�K&I��U��h�.����r��r'ǝ�_6���l��f��C����{$��dJ��d��h�xS�u͜Oφ��<��#ש^����l57����s;'�˾��)�|�$�ڇ��ӿ4�l��a����t`�v� �����!��,�%�A����s�5�Ý��N�k��i��ܩC�tm'@9F��|�����8�e�߲���?�D5sm�WiW�+�e�6ׇ���h.����k,�F��^V��l��~�����+����^�־��
�829�b�N�=�����,��E�ޅ��5&Q�k�kl��j�v4W��B��H&��,k�������:���Sl8)~�Q&X{>2�oU�V�L�_'���Vs��hc�\m���S�#z^�w�W���Vò�#mH-)e�֭m�\�5Z���g���X�}cқc�����L��k>}����ӂ�Z,���܎Q���yzI�4lsޒw��TR�aj*k��cC&�T9y�}F�p�3�v�,h��!88����n���n�ŉ�6�L��l�������n�ȎIɴ��۫Oʌ�gz�M^�� j@��$��2��]?���V�=s�蜣Q F��ͽ�y�4t�f�)7���H��x�D9^�VvOf�����;���	dI=�.��`�u� *o/S����mH�(��-(ұ"�_�櫧l�Ө˃���P=yT�YcWB����4��7`Ar���޹��B��G؄�y�R�*�O�R-6��*>��2۠�v�I2Pro�ڄ`��َY+�^/����j׍����a`���:����	1�3Z��|B�=���������Rұ,�&-�Q�)L\f��-}Hjg�������G�d�$Lku � 1��鐢1�G@�$w8�C��H��[D��jK���&V��8����M���O��;��qȇ���u���c���<3�F�-S���\�+�S
��ǉ:T.�>7P���:ý��try�ZbOQ��R�g�gK''�9�5���/�d���!n�8�*Z`f)�Y��N`�)� ����=Fl���y׼_�=��`3oad�>��r�{�t�1���J�=�̾l7�����q�6�gY"���`�`�#ဵ���\����$����W�^JJ	y�1Dؓ���&Wg,������Y.O�]�o�S2��1ǙYK�B�v�ǜn�Y�'�����16�p0p`̢�3�).�2K���}L;>������lR���kQ����Qs����˒r���nKv:�c�hRl,'mFZ6� ���;,cՅ�۸��rl'�m[WE)���ɀ{m6^�b�s����]�vŞZ��8iu��BT�suיv�������%��i�m��1��{�^0G�7_Tk�ԙ������B��ie�6�0���{������-���4`9k��w$KY�Jȭ�ùd�L2t���m�=�����[�Ӳpe(qq�y��g�#�Y@���2�B�h�Ӳ���u8�KV��WJMI��s���[8IO}������[T�4����':fW�+ ��rƷo�
c�}(i"�F<�6P��ө�>2~1��/�3�����Дc#`]
_��n���gi���ȾB��õ[�I>��8�b�
M�+~�����s���ZW:r��8"��R��ׁ0��ty�nI�u��|H�-����7��R��O׭7��{X-gm�U�{��HO�7��rb�
�$���h���4y$�V�g;��Sy��7#��#���<���1x/�W�g����e����N@m���};u�rf���zm�ʰ�>ڷJ�`qry��'ш{* ������]�Ͼ�ߝ2�ȹ��^t�Y��a�ש��u]q>��,K3�]�+����+N`@������S"��Sk��+b��&��EIf��qT{o�4 S�4�� ���=�L��T5?��M�ד:�b�%%/6^���'�}��3�˸������VUɈ}	�ú���#`ӲW�6h�������������G�wy��=�.2t푱˯�����fon{+���pvl��>��ecJ&(�W�Oa{n��Fu�ʈ��1@��hQ�-3���_�����7�0yKtMd�=p�k���������Lz�ӻ䎛t��]>Z��`�I����[^1@
�g����1�z�|�	$&��j�3h)��D��h�t���,ZcJ��
,�%��eW﷝���㶑��J4��"<�܌p�sj��͇�q� �p9?ƒ��h G���b��:*��9���sӞ{�?)r1��^��Fc6���9�H�f�����K��=�!��~]Klbm��3���n]}bg��Scll0������{6�=��3w"��R�#0l���3��]Ѳ	3�Y�K�:�yn����G��:�j�$4�~��c.%�ϱII���M�׹�<�Wg�<b��E�]��g�rnIu9���{��b��f֘~H�����3OU���@�6�$��\a��_�L�d�L 0@Ě;�xT��Ҙ���Y��k�R�"�]e�\��1�A�'R�{���9�ۘ"�����^��L>_N_
�@6_<6WIz�
G�*�
�8Z4�q)��p��@�q(Ϊj���"�{ՙR����ߪ���uo��9m1����y�&v^�L������{��մl;g�����gKO_����3P57�s9�j?෦�y�%�����k��6F�vsfT�t@(m2�3/����ԍFq������z4���H{��)��a�3ji��	���M��&�SӤnO�X����z��>ϧ3��[9��L49�����;����{�^��\.Mzr:��;��1ƛL��R>dj��D;9lk���m�) 嗵9�K
��^_�i�F�0#�mj��]�[�=5��1V� �	oj:?�d�4�/燈���L���R�D>B��ټ�h�P�R��2y�ԝ��NE?zI�/�Ϭp ��g��*��7�el汨e��m�8���Z�mQu�2��:5�C*'o�M��2�j�q�)�9H�c����f��I����R��?�xX]� ��t�Ʋ<��C�j��w��`�k�w�׍�i��tº�%���ܱ�d-�vEXܲ`q���ןʹ�Z���q��]�1�;�	������C@�^
��1C;A���f�:sD1��9cj#�9��;ym�Iey�ys3��ҙ����
����[�ե�Qc(S����΁��ܒ� `V-�Ǩ�H�_{�tƜ�9�t��ᢁe�`�F����x��������7�~o��gզ�mb��~_������cM�����FX���;�ϝ���J�JĎ{���}��ί�3r�OP�l�O �6�҃�Կ�w=��T�$�a#�4�1�����ǠV�o��������dv��Asخ�:�u�F��&ӹd#�g?Q�d;�[^��W������>�Mֻ�o�1�9�=���z�� S�)�h��?z��1;����c� '�n^s���Y���uͶ�3.2+��(u�[��K����
�dT [ת~����M�������ȟ��YY�fG���zY�M�ʑ&��G���1�ҡJ>��5/������9�׭s���Z,O���|�^4�+����7ckJ����t]��㲮W\���8�=���]{�Ed�i�+�u9�����̳�I>d�Ne��s�K���1����Ǹ	�.m�����a]#N��M�� d�-2���Ĕ�l�/߲�yr�!����3g@��]'�ܸ�&��.F0�9֘�h/��B�D�K+�aR踬g�h��־��K�f�)j�#�f���3�E�i��	���X��k�Ww�:z��ϱ@7�ߨl^/?�n�{PG�dڲ��������ˏSU��X(�G��=Pcf��)����ZG}h�!�/�n�\^�������R䦙_#�E��\" ���:��aZ?��~�| 5�ظ�PK�p3n�}�G��߿�s�;:���ڢ��G�i0fb�xyy�?�/�lzC�8�ψ1�۷�x}}Ms�sX�'�kR��,n����8�g�b�z��m�4��Nj;$�{S��O ���찂���5y�j�?�%]'��y���^��j2�~�����^n_���_;�K׮��8R�{ɣ��G��28|w`��X����)/���׍ʗ��d��F�W�d���=�v$������Ep�6�}�m��:�H��b��F}��1 ����m&g6�Z2�{�r[ʽ9X+���[�P	��s$Pm�O1HSƴۡ�Ʀo�Sh���]h�ϑcj�.��Xp�RB����&�AE��P���YƘ=�_�C>&��, �aܶ���;�bȐ�c�/40/s�yɌ $1FĐwD֦��������`o"�b����t>y������=�h{$��q�����������K��hOY�r��+{�M���uK�I�[֓?ә�ֶ#��o��=̖���}=R�m��E�6N��3�5�f�?�6"]�ir�>t˦����5(ip�u�,�_���n�'��϶V�O�d�2����=�f��F���t�N�|8�,�@���,�0��1��YVug0?��:HF6Qo]��������6�K���yI�{O�d�cN�ߴ�깺��#�Q,�&��ȝO�&}�<"���@
���Rr���uh�?k�q�>x9{L)����?���Zbt�Lk�3�L�̒�怿E����C������I���#�ZO��|D�:.����17���uM�^__q�����,2׵B�ɣ��B�#�1��5�}�*�ͽ,-p��gJ	u]�l!k�%nYp���a�l��bh5��|O�����o����˲o�t�HU�<ο�l��J8X����������#���K}��=��&��|��ϖ)Y�����#��L��#��n\�\�f�p���03�چ����N�N>t�ʙR��Bq����59h��k�OMz}�e�{2��W�w���40��6�G��w��� ��ijI8�����w%��5�V�X<�Y�c���64��gR��mX$�e9����;<�����	��>��L��f!}_Ľkk��u]���ϑ���2����H��9 �f��M�1��V_����|��x��d�ᲉkfM7,Wg�#��#�`�M�[�����k����Ǟ:�����zԁ��!��w��&���<�ɼwP��6��L��ő�U{4:9M�rr]R�zK���G2�{�<je���r����7����2Fiv�ދ��A꭛��1uG�Cv�3D�?(E�H.���!{���Q�>P���g	�O2I�q���_�>xx�Ν�+Sݣ��Ƙ��!��2%����nʛ�&�� ��hh��g��jS��ݾMf/�/�����m��Y[���G֓�.�o�f}Dl�ٶ��=��{��yF����>y��ɖ��Ӡ�-�=�,F�2���#�ﻗ�����E#zu� N:��s��K*K���X��%�"z<B��!-@�㐠��#o�fL����{/����B�@����K 9����x���CXSf�H�M�dk��[���d�={�@�(���4�R��Q1��c�'�=;.������lpf��O��� ��a���ޔ<TIO�7ʈ��p�`��B �6K�vTg<�̏f� <��{l�x��2ExK�6�{��}W����v�G�i��Zu-�o���dB�,�Þ��!���]lGϷwo�J��ߏ������)����<ET��%�ۙʞp�9����r�Kj��u��X�������ן�g�@�KL�i�°-Gs�6���@f�O9|��F�R�z-����/(�Tm*�ki&ػ^Bȓ$K�"��-u't{�"�%)߅qss��[��o	 Uʹ�p��bW�=��3�����g<J��<	P�;R�/��\?
�,Ai=��y����]P{�H�W�{zeζA3/��=�����o2|P�<ot۾qj�c�-�=�m���cl��>��2F���\J~Z_��^{�ׇM��H�R��>5��{���Dd�؍��h�U�5��+t����hsKǹ�H�#��H����y�<�=)��@�����M$�Z\�Q���<���6����l�1�!kNe�K�/�V���d ���C����-�r̺LA��% K���|J�9Ē����S0�3�;R�%ځ���CQ�y>�	J�`��i@�(�{=��. �>F}Iu�ɔ�'	jgD�������e�&�S�	��b?is>3q��J���&��G�f��G�9+!}!)m�gw����{��^�#�X��矑��B,7�{l;֦2�� G����{�����;T�,�{Tz�^ѣsz@v�Q �#�՚�:(���Z̔9�v�1�/r�]�4^|���͉4�8�1�뚲���?{�,K�{�ؒ���5'���ϢU��)@&  Z��d��d����1,��m�o�L�e2J9�傛�{�Qg�ĺ�U�u����2�㪳^;7�`UL���&E�#�J���uŒ�T�@��=�e�G��[���`f^���3����{�O��z��֘��j�8�?� ��{s>SHb.G�{��Bzu� ��<�� ��g�cV��Q��L}{��%�O�]N�o�Y�S��ߛ�v����[_H���^vRL��3ڻM�\!�	`y�$ �'£�?1���3w����1!��Q�e#��"�B�:0�7��Vˏa���f�5�������������{��^==�֕�)+��#����\.���R=�h�U�W�~�&mFf�MC��|�.ː�롺6�N=����}Q��;��L�9;oh�11�l�Z����cJ�9R����䔟e�/5�L;�w_���j�h�� �[�=˒����us���PԚ�R΍fX3�&�3c��J��)A
�w�9j�k2M���߲��`_�5٥�¯�tj~�79�|�I�ig?��	A���'�� YOԾ-y�)u���`�#��໢���o8-'�S56/����|�i9��PФ��.0�f���@�>8�IuB�rѺ�٘�Ӫ��( Z\Ξ�TI��a
�K��s�^^^���?���{��޽��؆q��޵ZY���)�����ʒ���������L�+��Uo��'g�t����v6c�=����9*��{�Α�}H���J4�ƍvކ�f���幣{�c�כӵ��=�HO���������u����[��e��J�����ʽ��v�����d>��<Z4��v�6��2�{��^�@�-��G�vk�bq�l;_ޞ�}��Q�rh������Э^�˲�k��y%�
�g��B}���G�ISkݲ5���Q��2��}�<�]�JP_�݋�6�F�����zqN�[�/m��,Z���7�N�fq��5y��[c~4��,i�H��Fn!h�l>G���uv�9[�3�ʣ�ǥ�~�}���o��u$U=퇦=�~��=�uM,��%%5��pf����O2�C�|�^g4kyǮ%�%����Z���i�р$�g��!մa��3^�Rf�� P���<�	���$��=�0.�\�|�:�������.�Ҟ5��g�y/9��&G�~^�ǩ�l��y�>Fg�M��uA�^���2ݤ����!֜�����ԴUdp��H�#�2�RzLh5�S�ka�F��|�'���ɡ�9;e?n���ZX%��G�ǅ0�!	Pm�<�SV���6�T���X2��Cuw�q�_��țvɡ��ʹe����\��6!�f���[ ��N%?ό��7!���M&�[uR�b���0!eg�Ɠ�6P�b��2jk�"m.�ھc�;���� �U�Ux�%Gd�V���ݜw���>�3���Q�e�)�<'�%�Q;�2��z��0�{2�Q�,笌�*�W�s���� ��ybME���5���K]�s�H��(�6��܂�%?{Z68�jBe(�>c/���E>dFc�A�@ҙ�كԱ`����`�SFf��PDk`�Ub�K\c��z-;�eI����_�|�1&u
k���
k�'7B��&�&�WaK�h	�|�����Rxe�un�X"W�S-�g�}P9���M�L��$��l�^E�w�]���j��=fp��򸚘��_@�0<�v�� hik$��[��ԏ��en���B��`T���� ���[X�Y�L�G�p��\<�7�'�S2�Z���2���f�����s�_���3��^��Hf���G3�Uۏ�U�̴���zAs/�gD(�:2b�\;�|��i��9#V�Kd�v/��ג:{�̫a;'W�cLL�`6'��-u5Z�Ę-k��t*�eo\.S��kR�_�k�/��u���f��gИp�8&�X~����:����n��&D�1	��8�]��k9�y�p�4��~�!����S��f��d����ڄgHe�ƀ���C��U8�:�.��K����c�c�Ar����=Bz �XcJ�O�}�����N{�Fۍ�utp��{?�Ύ����A�c���I-�%_Hx�1/C�p�\���F�[�)m���Gʨ�{~ʁ>�]�7D\��l����3�X�3����r$n&���~k���k�Iu^����3�|��4�>˺yD>d��Ű��@屉S�Qcr��m�rK�mR���-�D�Iz�[u�dL�
H�;�ur��h�͇;�鹤�o^g$���p�x�,��3}υ�Dn��e�%
�q\�'x��E�"'t}o5G:_$�T��֫������y��cŞ�j*4�v��=���G�H�!뼥�Q(�D�I�Q���=�Ѧ���P���w�gZ��/���1����l29p;�߼�Y�j�?M�w��{�/Ey�)�`�DaY\Q��Y�)�E�]w|�L4��K:��v�����|��<b+9
ia��Yleyd
��4�w����VU'�Ok�Lyo-�]��ޭ�ec��)�z�<��8��1��R^�G�d#�ܐ��}����
B�>#R���5*RR6��L��Jۯ�s�[M��[E�ی1 9;��)���Em�kb�9|��7L?�&������M��6�&����^���W�?ss�86����1L&iµ�- �d��wM�mgګ�4��91y�c,F�"��w��	��X�Y%-&�H�7����R*����E�Ci�2#3�d}���xn��lgg��`�gG��/}���-�V�-L�Ƃ�d���nmގm.��p�pֆlT�S_� ;6�ԏ��h,~[nˀ�r%����Q����l~f���k� ��UZ��h��+l��ţ�H��~�ט�=����cqg�<5��:/��۾�>�Kft��L�G#Rd*H>N��]��5��8�>~4f:[�jȧ�C���t�����\S��ybm��cl�Rr֘����!�)��G��I�8���h��S�:�����0��@Rˡ\:�����üo���r��LV?N�I��fh�����Q�ܳ������Ly�-���s�*��sk}mlW���f��ˏ��
�h:���o[�='/t
aHc��$��l��o�\7�c�\��G��<BB�wko }~�O�j��薥n�W_t�vj�PC�.ha����M^j߽6�g2���\�,K��s����0��k8~��! ��-��ײ�Y��L*k�*>j�!�1�9�VY��3xl'��d�)ؓXm�k�m����[U�#驕�كd�~�ro�ia���7�!�}ɷ�����)�2��>���
�r��򈴬������)<���o)�$A�������u��ZlbY���_Zg��:��0Ɩ�;3m��T��A҄J����5d��� ��kOz���A�-�m�[���'3i~R����8?��l��E8�Σ�/����
gnZ#����e��H���y���S0�C�.��x�y��f�cK�%�%N6{��8X#&zO��m����-���{.b��x�E�QLZm�X%.7qsm��
d`����b(�.R�I�T��=%��7�g9���Y�����g_��f b�+�����4K��m�5�K�6<N��me�))Gc4Kr�=���Y�ʘ�#���ïkQ���)�Q5��������t�A�A���_֯��40�嗒cK�ܑ"`b�E�>/^���2Ƙ<ե��I�0g�L����b�C��hm"����Y?DKk&�U���:�k��́ʙ��|�j��A^�0�����@̡�F�Q0��菪AG r���}��j�0ƨ��5��s!b���b�-Sv��W^/��Q���8��mH���'�X��Fcgo"�w[2
��J��m�طv��bv�i�����=9��炙�����Z�ey�#E��zA���=@#�9�|DOZ�M�<M+$7��:��t^v�3Q����w�5�B.���{�1��DL����9XkBr�[��6�14m��;R] �����x}}ů~��]&���Y�C��ʇ����dd�+��t����I�nrw*BD0	,Ri�%]n!�ؗ(��f2�D�T��,3�@�N�v�r��-�IO�����%��v�-Ձ���|���Ytf�������yKn�{���Z�hs�Q"mB)k��E8,�,�~��Ə��#����^Zm����6��Q�̑&`3���ϗd�����h#b�pnA�fcy���$�����1F��o<����-��'m����|LƟC��r��iIQ��k(/��M�������:�0�$oc4����[vCs�8"�8�h�]iO-1��"*��G�B�G�ނ�cb%}G�z�g���`��wi+��3�s�v�.�y�����-���#�/��K�{�G��#���r�1��چ[�F��ZM�L�$���h���2�:� �����qj{�>�e��/�+a�u�	�d��\o*�2�{83)������E����! �l7�I6�н�rb�)���B^f��d�Hՙ���)X�Z���pʳ�EԘ����cw���Y{�{�����q��zk`����c^n�������ɶ���⾒��<I�����p&p���P��÷n_oӡ�x�u3�r�~߃��գ�����{V*�!�Ć� FF4��ݮU�k"��� ����{��$�F5���e3����a2}(�҇��_��q4@���Te��j�Lz���L)t:k��dOQˍ�^��]�s��u�p��|N�x�7E���s)V�ɞ��~H���Ud�k:���JH���	��6Ȳz�^]{����
`���aO���}ǘ�=�&m��G
m"�6~�s�,x=б�p�so�2���Im��3��;Ƞ=��6��l~�ؑ�8V=�}�MGk�nFn}V3����y���B��ݐyG=ӭ���9K�OH���،4�8��^���q�O�0�9���u-ߗel,9�-�0��uD�6���~.�a���{�~�_}���u��Rϝ@��%�T�{�s��=֐��?,��	�S�%�,)�䲸����b�wJ��J�]����w���Ҕ;@m�*!��{��G�{�]�6�֜���o'�=�w����ͤ��f���7�o��S?ocY�>�P/��T����cQgd>9�i�{����6��Y6sR��j�)�n�Gd�Ѳ�e&�ch7�V�[��2��a�˥H���m����S̮�k�N����'	���Il�dVU�� �E�����'5n/����7i�c{�v�W����:���^�&��{��FL�#ο�-��т>��:8�,�l?�ϷN���[OV��e!�/Ն=G������ݘ�|y���C�F-.�{>÷�wF�,���#�y���>���m��MEڐ�Ȉ��F[S����Wc�)BA���;�m�W>��\��%���JX"��BT�H��wOb�9�Fv�0�iyI)$MJ!I����$���o�iO9b2���a��V����3v1��������-���һ�+�b{ &@ٿ�B�F��d�-�\p^.G�M��М�M���B�v=�-��z�"�7_�LV���@NךԺ{�V�:�1��� �v�#�����ݕ{���|CԳi���^ �7ne>#R�3jב�z�W�d�|�!{0�N�	(K(&e�����ԗ[�1�����1=+)|�yn�����ڳ>ҧ���=�����`R̵��b���+~`�cL��-lcz�RM�ŝ��έX�����@%��Ͱ����_q]W|9�R�'�ksj�̀�k��"�A�3(ԇОGYFq����ba,��b�4j1;{��6��ߜ��_^^  ���0����e���A����R�%�����t�$_�ib��~8��2ơ|t��壞+�x�
�݋q�7$�5=���Q�nϓ�����`�m�k��#��u��va����a�&���>{e���v���H��|}��_��;k���D;�Vژf�ܼi��6��u{s�|.���7���#��Oi�����u�89c]פY�mh�G��ƴ����+��kW��s="�8 	�a9�"�����$��ǩ,�n"�Ӳ�z���alL���g����^�j��Kk��l���1&;QkG���+��'�x��hjZ�h�K�ֿ]@d�.�����pRg�Yx���x��9��!��O�Q]��ٓڞ���>�#n�r���/���t;�E�^�2X��c��#�%E� <ji ��	��󹪧Ҥ���Q����O�j��� ➶̵A���k���F�a�Z���Z�4x_6IG��y1�tfQC������M�#�laG���cf����h#6�_2�{��#s�L�H5�RX�Nd����;g���-ͯu}��$m��I�R�nb�;*ᢽ�&*������>[��c��	�k���֨Ww!=B؍��s�����[���&��:��6o������9g˿���ـ�$k��`���V�E�N�2��[ط��E��eE��wD4u=Y�v�6&����6j2S�U��eY�)M���h>B��S�˿%����i�zy��Z�z��H�ӛ�%��G�<���zd�=F��>V���~o��̈���7S�� h@�v���~"i��R���˓ą�)�^(�jo��<���35bs�5��@N#�O���!$�@Z���+�%���Z�2��c���#������pa5GY��Ҫ���$�J��\�~�PG��a�U�N�z�+��Ţ�%[�Ӡ�̃1F�hZz���>�Nk����T5��6|/cVu��l��F�I����gS����Y0�~��#"�����GJ�Q����
���.71V-������/���
h�t�iY�X�FQ[����Kf���=��sZ�{2��aǈU��<ͧ������K�xg��A�Ƙ\-�CMڶ'�����=��H����z؈�֖a�;��9~��i@��sy� �bbZ$M�G���q�`�NIU�6*�ja�Iu���,{��Ђ�<��)KQ��|릧��{{�����]�,3�k1����s&B�Ij��)�mL�m6�y�G���c�N�v����B�� �k&O����l�HJ�_� #��x�Ͻx�{�m7���@�)��2��[�g��=�q{l����s���h���V3�}�m��BZm�N��7OqBa�^i£�g���>3��&F��
�d�N	^f�Wڜ��1�m�H ����C����&(|�k))�:ޘz�4sH:o~��}��t��Z�o߾�z�¹?�����;�iYpuմ�r��q:�p^�~��<B�%��1��v�H�QY�~�DX%�>�F��@f8�m��f�a�����0��v�H��5��G��}�H@XS��l2�6�4 DE�.U�U&��d0��ϵ��A�̂l�v�U�4���hg�s�h}!x�h�g<�:6"�U/o��+I�[d�0G>Y'@�z'P��n�@�ilkAߩ=�oΙc{RA����k�}_�rt� m4v{@��{�Zb�s�P��^�n1�l�i �f��ic 4�T�kڱ�3�u6��w�s۶[k���1)sac���e���QN�T�="'c�����c��5J8�D/?x�҄r�!c��@R���_a��.g�	gܦ�'\�Ks9
�nW�6M3e˿o-G���g&-7�l2�������� ����Ԟ7��T�g�X74�S�H�צ�w��>�KU�( 7#R�XƺۏM
(�	;��Q(65;ͤ������|�ܴ����y6iv^���#uͳ�4�;�����L�c�~�"���������=v8�^&����#'_M�����,�]���BV9�R��`���XI�7��7م���xV큵����6<�d&�cm�����@�s�:��HJ�t:����҄;�]�'=�Z��I�4.�����kO���H��N������ˏ�s�|�ލ�^�O�kpZ�ͻ	1�Djݎ�io�j�v7�=}?{f�(�:�eN�J��1��7�x�O۪��=�f�n�BcN��
@eI�l�gC7im�b��gph��Z��)��c�3J��8�̴{o��j͎�3�G��K�W%�I��豗�6���z ��!��H ���iS����eLf2�3��N�VF]g�+ �{��x�Ǌ�.����r���b,L�@0�eA����\8�c�C���Dd �,b>����ю>�F[�:a'F�Z����eO(��}P��/��kvp�N<f�8�B%Cl�S� ���i`r���57���l��.@q�:�O�{��@��}�=_�9�8�Ok�d-fm�o����S2bc�(�+Q�+
�4w�Tm��yΊ���Ҩ�ӱ�Â6�pp�x�z����Os����coCc���(v��S3>ՠ����w��������0/cV��t�������r:.��r���5�l�0	e����W\.x�q.!��Ic�?�8�ۯءku����:�!q�d&��x}}�u�8�����?����4Ⱥ
s�����3n�>��'��$��h�u}F�.F�T�k�om
�.^�5�q��Sp�G�6q��"n�I�=��xX�c�̫�I=B;��NKjfJ�^��Q̝�u��>j>���݌�1�؉�]`��nM�J�`�7���������j/�\�;�`ZL=oiӵ��`�Ie��[��'�.������n���x/�K9.7�>��
�,^^^
��H���ܐ6A䤎O�d@{c,�Q��� � �ކᳩ�!2��P��d'�q�"^�uL&�'/rcڸ_� ��k��k���-�{>���X�Y�z�� 7��`�C�^�Iʣ݆� ��6eg��^��x)�K��#�m���HFuI�P�ǘ�;�
~�Ů��z��s�������{�㳹�����C�N�%1)"D�)-m�	������7�\�aڵ�zqg�l�hP�QMR��։ldZ#�-���ڛf.65�9�����xW��8�V_�f��{�B�bAϑ{};gw�M��Н��9�@'�r���rm~�F�Q�!�
p6�޷
�I�:�u��˲ Z�,�E9�:؎{v�%����Р��^j-RT/�� -K,@V�[��j��O���8�Ga�}o^��@L�����G���D�)�sh/ܟ����g�3��z���1r27���I��e��@M<J��>�T����z�sҽ �p}|�{���q���$kVT�&֤ \�H*���Bs��2�4i Y��깭}��ןC-�˝�c��\�qZS�d2�Al��31>���Qw5�;�$#��79�G�@\��[JG��C&� ��|>[>rΑvkj�b+"l�ٚ�m��#�$�� �\hW����Ѥ�Qf/8m8:��i�!g�=�#�^�������]��X\ʿ�,)�+W��}��g�m������q搳��)�c#xK������5�ܲ�	V���L��mƣ"mRe9��LǶa���a�l|xT۴{ؾGo���e��t�����mjYJ9�j���`4�������Mٞ�{k_ݳ��u���	7��Q�&�%F�b�f���V�y�k�oT�X犙���-^�ӂ�W��L��Z����1�@HF������������7��Q>ȼUF��O����;"�I;�1>�dӐ����Wd(v�48�%�^k��7���˺f&R�Q�=2��нs��ٲ�R���s�����V���hq Iu�f�dy���X����0t�#�hƾ�����秙��'/�ῷh��g�=U�6��L���f�U�c��}�bC���r�;���d~I��oo�)��15�>�c���h�k��v��J�����E�63���Z=?�b�}��v϶�^Ռ�A�O�C>Zf����,[�fծ{�磙�#ҳ�{Hٝ~����2|�i��~�&�(H��0��;��g+�l~�mS?%�`Ž�U�^w<=:м&2$�1G=��D����#$;�޹���U�c��� %6�Y����[�Z�0<��Yl!$d����fE+�2#(���k���]>&���s���Gm$���.H����ܓ4qP8��l�4�ײt �m&���utu@��C,񀲒Y�*9��<�\�r�y�E��ѥ��26�������Ī|�E��(K�6of:�����*c�U�	�%y�(�W�/3I��J|G݌��BP��h�yef^���3W=���]/��Hb���E�=�,�s����a"�a�۔�T�������l�[���,��7��[��x��d���%G�7!�L�t)�VT6�&[m Gk�|:�S����m��r���!��a9�gb0�9C-�e%eZ9�8�T��Fcj4�Dc0{��)TD���vh�1�)�O1F8��r��(�A�-�A���z��I�V9��Q��tw����QWd�=���\�1��g�j����|�!�)gL��Hw�����wK��X� ��{�U�Um&ift������8z
=�<J��d&�4mRK��3�Օ�{�� �X������q�r����$ ����?�1��Rm��ܳL� ��1G�kv��Y��wm9�8(��H�m��k[Z�o�ʺ�����.���t���f'8�vJ���2?�D���c�������b�9�����Y�m�|��A>���;��eI9��C���6�9�n7<J��P޽��mU��i��6F�>c0?��چ�b�~�6��Ř��%� �0x ��h�Ѝ.p<�&2�c]�mL`�U`ak09��X��3��dJoty�_�cK�|�[s�1&��z��A����h�w���*b�!{P�8���g�x���Žz��@�>��jR(�qY#ؽ�`��D(����\n�w_-��� �-3�3��$@���ո?�|yDZ*�3�V̺[���BJ���|�� &N�a���M')s��0?�2�� �"��i��}���T���E$o�{v#W�%��B���u)��4G��M���K��d^V��"#mcuVn?6ە�J�����h1;�!x lO���gm>��� �5��k>�8X��&MB��v5� ���Y��TL��EFR4�=��ۆ��Sq�*�&�.�䡎p}����WF�%��eYk����^[}�JMp��c�e=��8�WH˴��w�o�d�M��8��3���${Ŕ��6%��e���S�*k`ru��ԯ����ŋ�V�3u�Ed^|||t��������GU��0�@�^�F���H��6��{&4PK��<X���v��X���Y=ԯ��wK�&s�f�E�/͉�l��34MN��/?o9������ ���4�$־��h�J}B{��^�)�1�T��H����ʈ9Ǒ���<c�����aY����.��B-��~7����L�_t�M�䱙)�8��$���e��v�d��l:y��p%#�����o�l�"[.kt['���s4@aϋZ,��g&s��ܫ�U ��z�F�U�޸f��4u�����:戌z?�0*�Lrl2� qM#���6lL;�Z�-�*�3�:��9���^&��LǸF^8bc9"�򜵈�(`��;���+�����蝾:<Q�[��}�_#?#�g��ڲ<Z�6�F�֏>o˦��H��Ln��*OK�h�)�&�>�>)BJ�a��E�3��+Ь�]_r��i�m��>�=¼T����Z	��6�DՌ�t�p��/7��R~Lf�Q?��Ę:vbehl)���5mક��������!m2�]�����)�+�w�������{
�E8
������^���rl��r���Y�[�U��5�^f��m�{���᫄k*�z�0D�';��{��C���kd�r5Д��	ώEK�`\*�#�?�#מ�Y߸(g�Z��_%(:��=W���d�{�~�hy�<äZc�0#Y��GBrQ�sk���������>0@7v�	h��wV��dc`��TT-
�*q$��5E�o9�ĐlD,�isiK�ro{�S;ߕ:PK)E�{'ڑ�4�l5��+�LY=�~]��L�Enߥ�="�C�[)&&I�v��1{��}����+��I�C�1��,"�+O���9������u�tfo~DxV��*��.US��i�Ɉ�Q��f#��<�5��%�7����$|�=��U�ˁf�p�jJ�0���f/�/�\J�j��%�K�~� :
��0�β6|�pe߂�|����������&��`m
���J	�E��@����1����Jgb]��=8-�ju�3usVSͽ��e9�1����љ��˂j�oBǨ�F�!�+�^n+M���Z]j�j�)��l��c����u&�/~�����˵�ǟ�w8=;o��Y^�R����f��M(�F;�����A�?z׏��~r&�P�µy��V0֭u_Ư^�_����m	 ��%5�ߎ:�ny�k64 rE���k*�}�zH�	�dڕ�4���Z�T}�/쌵�͞r�\�{�@���Gg-|4�K*'��h`��p�--u�H(!�7W���&�XN5���� �Ѯk�i�:��Z���t�q�p��vB�ڧ��h�o���Ũ[�vՀ���Bd\Ŗ��H�DYwύ�{`%���@��C�n�����3g��=��^�����?K��~	�H�P6� �%6��ҡ��縮<���֋���%5��/I��}0C=����[���b4N�\���|¦O�v���o����a����gn�V�϶ ���n�|������0
�"J���k�8)���N���&�Ɵ?�uK<CVm�ф��Qy��MY&�����5)ʍ	�8�6��>~���ǌ�?�\�/�:}�w��2��K!V�"0�)CmPБ�4 2��ˮ��<���@�2��>�h��&��x����[��1� ��1��e��g7iS�T�Ҭ�Ȇ�7د���"�Q���8?�Xc���~=kà�H�H����{Ҳ�n�1$g��#|U�@"�܊��փOyY�b��^��ssT��m��`A*������&EH��&T��kȟ#}c�_����f*Z }n"�
��x�=[�32������V85~��^����P�Bn�W��Y���cr\(���W���]�Ee�3S��-kmz�J v)�y%[���iA�~��|R������ZV�1�jp�:��5k��oDk{iB�}9R�3�Ք{��i���N	�>H/{F�#v�Wm�N�)9�p��c	\\N�O�Xr����cא�U/��(S�c�ͫ,��Wއ��.ƀg���i��8�1������L<0~XxV��Y���2�����\��q��֦'%�M��F�#Z����� c*�Y�$����@6���b"�Ep^��!��m�~�*������"Pآ%��^/�c2cV��>m����A��W�ĘQ5;��ti#Zm������]2���I4��L��MenվK��S�W�A̕��M����L)dk��3`X:�h�k��A�rߞ�s0�Ȟ�C+KW�3bK�r�m��{��:g�2�z!L��V�4b�|U�i���8Hi�r����f����WH��>"�XXg
BH�btM��e��P_ӁDK�x�.͑�w���M�ga�DB��{<|||$3�`C�97�k�d�z�>�'o��l��&���$�Q��j���eY�t��v�1��	�Ӳ�3�T/)ƈy��x<���s?
m~�;P�T�Qa�
��`�g�;]Ȳ��I6v���%-���m,˫'ʞg�:�Z��X�^f.��*�g{^�g����e#uƃ����o* ���P�[�	��b���W�eU�<�� Z�i./�q�9_�v�-3��*��P�q����Ԟ�*�D�7���L,{�܏2��0��-v�M�ۓ�9BYw�=�_�i4�f�B;Q��^@�wm&0�E�m6є\������ϱ��ÿ��o�8�߷��:�=&{����k�C�E1W��Drs'2�i�E
�Xˆg�C��H�o����ͥpJ�4��z�a��W��x��Ƅoɖܣ� �PLM\�Ni}�9��P��~n�g��2ai���M�ܤFʓ�^�֣��w�Ȃ9V��U.��wX��w�N��Xn�����c��p��밒Z�&!��s
I��9��7G����1���T��X	�H����o,�����Mڎ��B�2���D��*e�l��vkq.u`���'�&Z�����a��!��5�#,�u	X�r9[�f���ž����;�I/s�.�� }��2�֞ﺷ��n@&�`p$d6s=9�kl�-���]�aS$��m���z`�\/'�d�z-�z�~�J�&��8�-�'㞭ɫ����\�ψ�l��3��d�ej�P�������Ĉ��l��U;�A�cs�b+IL��Q�g�Ej��d�z�ڷ�E� [�٫�Ei��'�x/��`��x���G�����
���B�u��E�vH&�Z�G嬚���i��"�Ŵ֔��˲��1�~z�pG�<�>���[@�Q��h`�Ê�&�`���X;��F�������b]@�K�WL�u�iO�j��Ư r��i��9��Iu�Q&�k���H[ d��Ԙ����Km^���\��'�j��t�s���ڢ}�
�r��N�o�Vi�)� �lf;��/2CR�0��D��o��3A#,ti�S\��3�9GdWU[������lëy=ke���/���`8&���f+�K�nƵ��f��V��h-�\��Q��W
w��+����(v��k�i`X�m6ׅ�-��n]��F
!P�'����'~S��=m�MZ��N��g�օz���1�l�0r0֛���O���tS������ؒ�Q4n6�A�t/%��4���i�2�|�E�9�Vc�Nc�@��)�?G�Ѳ-b�����N�SP�Ȳq�ŀY�5�;�z��]'�9]O��+��R��f�3Ce���d{���[���=\>W�1P{Zb
-5��Ư_�W��~/4�w���ל�r��/��V�!M8S�́=��eS�[;[m�9�[`��ֳh{���a�.;Ҹ"��{k� �ʹors��.ڠrV�	�D��!�b�Z�0#�dT��q�c�)W��&�['��4�Mnr�&3��eY��}������LZ�"69;�!(���JmkAq-#P^�s�4�ESQ��p�SH�8 ��Ţ"��1������r�˒C8[}��-9��hMx~ҫ�}U�?�q&� Z�I��doCj �+���g��8�f����u`R���>�U�G���-���rϡ&�/���,#'es���w����#��(�;���#�JΚ����iT�s�i%,�a���R[�w0?����.O��ܬ��-�`��Nm���4m���1;I�u�w�$)(ui$E��ï��l�����/�6�;ȷ�����]c-K��#����V�g�drN����S��-[����+�O�m��W]ޓ�Y��=�,������B�� ����=�	�L�nU�լGu/���S�sYWP�����Pô�3G�Jq!���zr���e��g����w����$cʹ�[La�Y��~�W�% �l�w��uZ�4E�H�8P�1���9;�X8\�B��M/�L7�ٴ.��t�	�W��@�Վ2�Z�7����,��{,�cY<&_�^��q5 �`����$�~.��J�2��W��R].��;�Z���=�T	B��fl�]���ՠM]EXǌ����ᬪ�/%U�1�nx�^?g8��;H��T��D�V��oi��g$�`vO���A���n�C��[FZ��m��C�W��#S;�[��I��dd�����>��uy��!�6��HG�>����Vi|O�a����^vF��d�pa�Ċ'�5v}���f�0ݝ򌦗Lq8�j���F���Z��B*v�zJK))O�������m�0Z^�5w��myV��a�:4U��Gڨ�������Z��7���nXPIF��=P� �*�v��f�xUg)�b�o�8R'0�!���@S�K�d�m{(�,`�+݊����1g�o�1�J�F�)`��5��S�!��e�9�����P���T�k���l�XWmf}"�}�5�T��������!�F�ԍ��v}o��ep#bD~��{,��;��g*�烚$Ad�_�~^�_��`�?!`�&8����w��ƈ�Ci�&��˜�g��X|�B*��:�4%�l�Φ7#��'�^"oG�����廯�� �L�9}���z�H�u>���7�j0���s^!{6vWd�9*��OڙY��V�*�8����Hf��-�;�6OڍJv�_{�ܯ�������3�\�x�M���?'��N%4��p����$=';\�L�~oB���ԋ��~��"��l�C0&�dN1"�m �����3��@��c&��PK���eZ�w�Ó�ǟRƽ��1̀�hv	Ƥ�#L�h���r��k��x����O���UO\)_�`Rl��ܳ�ܪ�%���R�6��h4V�hF����LuLȆ-��sa�~5ֆ��G��(��i��ϓs��5����H{�����ri�Q��Q齇V�̞<�T�_�8r�pJ�6`{�ܓ��Pz��k���`w~DF��-��Z�Ϋ��T�5����bnI�
D����~I��&���v��]�XY" N��M���+@gK6���C�TP�X�Uv�=9��&^��a�u�N.��qU����Ssxfc�"zB��e�_�����}G���["��˟��oJ; Z��]��o�o��*�R��o������+��J��.�Z�j�Q�s�@��9�=�1�98: ,��+U��5�z�I�r��R�61�^d;7��<g��
y�i>�-�!���1�� ����1&@���s������)#�c5Ho�[)�r��܄{������?�v� ���lr�B#7w�1`C�w=aI{M�Gl=��xy�E����j�i�ک����j�л*�R�>S��5���|&=��ݙ��e9�mi�U�Ā{�P<�L�s��H� �|#q�h��vܩ7	�.[�^����'��)�i�v (��˩lelFR�O��Y�ϝ�r��o�m�P�s���ٰGbn��"�X��&������M�G�v�Y�2�ׯ���lG�)gm4�2V��h{�|z��(<k-~��7|~~��zŌ�mMe��bjgMq���8  �d�cļ,���X��V�d�����H!�k�����L����`����K^�9�Ӻ�#�K6a��5|�N�Od6��|F��՛g�c*B�T�ʅܽhjI�X�'���x+�u�
��r��i�P�_��Մ�Fq�R$��ǂ���B���K��lH���^�s��ޙjO�&�]�m8��(G�t8�Zm�Ur��2�I ��٬����	���&�%�f&�
�$%�[(sy�ޚ,����o��</E�-�=-a]�t%=��w�ny�M��&��=���r/�:5���5c��L��ck�sFu+3���Q��_?���+s$�c _4z�����i+,ޞ=�Z��Lk��o��E~nh0�TY���)��6Ί-g׮�v�A���Gw���˗2��u����Hg����˓�e�N4�ƙ�7U�QVv#�;Tc#�E��=�Ɉ��q�������h�����_!\[2j��/�j]�1쵩h�2�Qk��~����_1S8���#�f��n]���B�g����n�)��w���d�|I��� �(���N���������ZГ#������Q���0xPJ;�V�3� 5��U���:
�Yc����P�Y�#�7;-V�+���k	�e4�W��oL\$�Ǣ��5���<??lK5oi���3�e��j),!���#lҕc��+������s�d��)u�5�,˂{ν�{o~����"�Z�� Zz}@��;B<�М�݆������A&7�=k��if�����a��z�i&��Z�©�PT�6F h���J�_Yw��M��L�iN��rm�u��5�-T;ZY���lSO�°w���q�֬r�i18G�15���"W��94�V�L��~�o�o������}' 5{�L#���v-�e-;�	蔭��g��ʭN�\��1e�m,��ʳm���K�1y�:r����%`D��%�C����
p8 �4ֿ�O���Kx0��ؓݦ�ZR:4�1�����`�{�0�w�'���!�`B}[���9JD||| _���x�<R�k�"MYʽ�? ���c���2�5�Ai3�>�\	���8L�����>"��<'���l�a~��p��_-o����|Oȹ��
x�̈́s��-����/Y����u�Ҍ2�����q���)��?fwt��9��]Δ/E2�|�J��f�WY��C���͑�+�
��y+M�T=��>����H�<@έth�%�yH1���{v��n�dsN>���?���Z;��W��!%�Q�Ǖ�O�� ������ X#� �P@�|��.f泬�^*\���Y���|_�����೓�4MU:M)5q��{yd|P��\�솯�2�����*����
.���<g��=�ɷ ��:T�����G�Y���W��D���E�e�-Ϟ��'�d���_~�ڴw��ZJ�VmÚ~]�H����l.-9�QZڄ/�Y�>�0eOf�iټ����Տe�#�z&�^�����AS�� �̐�Å�� ��3�)�;�,���o��S-ryf�]�q[o��{QH�҈�U���(iy���k135��:���1D�]i���y7�7��}V\^�)�$%a�h<Y[�HZs�� 6�!=ᚢPއ*��V�fф0�,���l�A>���1�~}�Ҟ|��?ϸ�s�nLbL��@��IV�'D	��T�2P�Q�ML���n��6!�Hk ;F��a�5�N�#��U%`�
�63�t6�gaS��r�M���
��MmA�������d�E����1$;G�)�;b�"4hk1���>��k�u�n'��f	p˾��}@:Gf�__�a.ץ�u�v�z��k�5� �Y9������Ù.�.m�+ ��xv~�q=ʨ�LF�0��N^��i�k�e��Y1֔�4��4��g:5�^ש�Y�� M�_�� 0�� L�Jk�/�7��L�=���T�]~Y��1�?��b'�N+�<�r}���Z��cZq�V5f���<�<n �������f���7S�|�6;:��V%�톘��>=m�¶ڴ��Y��\�cȭ��?�=.���|�9b�V�:�3�����&I�j HdU>s���׮8� @�X������v�T��t��7R���݇����pT��]���y�M�..�CYlo�G��}��	�k����( \9�J�v�N�@e[����.�E���z�(v�v�pu�~��j�D���Fڠv����6�*�c6�π��֪K~�.G�՞)�).G��y�S<c�����V(�������S�t�֡��������}�C�Z���矇���[0��ך�C�ݒ�$�t�</�u�5n-�e��mRmx��l�k��g����:M7�نK.��I���d^�Jm�-� eqƦ�n��m�@��yFZሎ�ؑ{z��zX�01��n���>������ل��� [>#F,l�k���T'VNE��bDd=��
�i}�I�Rw�HƗ��8�̡��^�=�Z#~���VV���Fd��_����B`��C�����&�>�\C�yzb�mf�A���b�^͠~��d�R�;�tc�.2�,��48.k����r�[犇�W��:l��D*�d������`=�gge��Z}n
H$�`��j�Q� WN��xiq���*{�QB
1s���lt���'T.=O�Q	 ��Z���ff���3��6�{�ٖ����sf�Z��E0��0v�A��a��}q��8�դ�5q�z�jeI�V}��9*�/���:�R�����ejG�~�{�����7�=��}���w�3m|v��s�٭)�Ѳ�s�ޗ$-n����y����U]��8r�=�w�o�����H��(��|����vT�5K�x�Sl�#Z�d�y�>���º�Li�wV��ǁ����b{�6(�U�&�C	4bV�l; ��&�9P����ݨ����f�f��
X��9c�^�:�{�S��CƙQ�1�WlDTƤ8d�6ly����Ze�d��5$Op��jf5R�]>���BIS0
BZaq�������K6��:�%W�_����$!��U}��1S���{�	2��ۃLm��-Ĉi��MN_�6'����o���7M�,��a�6gL��4�Ի'#�5-����[D4{����8�i*r���՗�����li3��`!�+9i��C���b?���d	�g�	4��m�I��'e�;w��^�}d�У_�S:���-�ͳ��g�������s6��S$U�d+*�j�����\:�w�k�Q0'�.b�[�����w�m��{��VK+�C8d���-�:��@9�����ڒ���&[�V���m����)��Y�諾�a�x�P�[ǣ������v��=1��wl��V���)"F_���r&���(����}�_ҴfO��V�K�=��>!��*�;Imd�@�Ń�;;\Z�P�92_=�j�a����m>���G��U���,t<�n/���(n&�<��V���  �I*r�Rywyo-����Py��pDPHfJ3��'$&3[2p9wJ�N -ٲئ�	��l7y���|�X ��U�ً���g��S�Mٷ�һ���rj�?69�l��PS
a ��d<j�5��1�%.趬-� �黳]�b�FL4�v2�A�w���ײ��7��mAffU��ggS<�r��u��ֹ�`����G��B@'Qc��0�S#'���[6-���(��듻��-U�glr^�T�=��dY��2�%P;
��ݱi-�+ ��+ve�N�mB��!xL�Y�+�3�x�v��"Pz�@ l��j�W��{��f��L�Hg�����ڃ��H4�{t���i��@s���Z_����4��d���Z��l�w ��n�as���ĉd3W�f�<��^�J�����G��!�����i�Z�	���{��B��{�i m �m��Hu�O۽k{!��h,	w*ן�~���U�}$�M�-��1f�������Q�i9m�6q\=����F+������b�853o��'��6���h ���PS�6H���xm�{g��rh�c=˿n��2|�Y�}�U���Je�C��c{oR�r��?7Q5'�L��q2�5<��=�7�2i�]C�-o�6��GD -$�&�#����B�`Z�`���b�"�I�4\҄-/Ś�^R_����u^nk�I��3�΍��c�Xj'h�N���rn?c�g��-`�c$�߷!���F���zzR���l3|A]�1�'X���u"��.��(�3�U�U��Q�pL�i�ש>c�1f�ݳ،�wj��=��5��2 ��:{<9��Y������7bCX}�h���p�q���F���ඪ�m(^��ًH�s�.mȩ���%)e�����m�is�`Q�Ǯ78\74Q�� 6�G� a;��V�
Z��%&�m�&�.�����Gs�k�ǔ��u�Y��-������ZNc��5�L�/�DRE��.ʫ�忝����U�l)i���������o�����C���N�&L&6��3wX��t���'�}�w�W�ƯTsH#���s���YA�Z���ǳl#�7�!�Q�fމ9"�p��.4�e�U�c�x�9�Ԫ�P�������RFXɖ��cm�*�
�����s�fM -@ҿϻ���=S� ��{��e�t�*kWc�msO�=��*;�+D:M�[�%�ge������j�LG��%�lfo?�x�Y-�\'���C�>�̓��֌?nr9����d�	g������he�S��k]�'��:G�c�S����ȃ-���L�=���8o {��P�
�w5���0J���vރ���3�{�#���@�:rY24Shj�1�r�vn��sа�	�cfI���jcn/���8%��y�Ҙ�hOQ�✚[�J���ς��7!�k4���>^�t�6���3�R�O�����I�"���{D�4�����ޓM<ӌ�P9!q'��w� L�w2��f�����y���?�F�*�p+=���="�~MS��ޅ��jV�l7� �BQԛQ���`p��%��ۭkG��8�T�G��9$�k�[�s\Kzl,�Wιj#k�y���Ҳ���l���}�p];��a���]e���ע{��]����'�:b����8�Wȳ�Ƕ-e��8I6�%��ac���}����IZ�6�~���<�/�K�Ý���LkR`�^Bw-l\m)���3L�`��7�4�p�<�jՅ8����)���jK.��=3���Q6� ��#6�����o�쎴��3qM %KHK$�I�m�A�BcO�%g2�T,��N>v����N�^-wp�p�l?�* ��Џ
���@QS��يg�;�T�ձ���[���L�@��3���Z�n6Yze��s?؞��
}D������#���ޅPL�$��BQm�ֱ���sO�ѹHk�e٧ �pX����n���� �L5<�l���ԥ:~O��|l��sA�#5���&�0�j��۷ۄ��G�,c������W���y�1-��1e��4Mp�U1N�i۬���%��Y�x��/�d�dc�/1Tݨ}�1��aU֓E6���^r�6ޭ�^�����W��l�3��"YCn�I�gO���$xj�QG�Ƒ/��H"Ǖ��-�T����6�{"�Ƥ8?�\?���K��gee�.p����GB���?R��Q�3mѼ��FΙ:-V�l��m���7� 9�*7�82�����lK[��(s7J4�B6�O�����j�a���]Il-˜��d|���u�`��?��0M�M���RP��5�m�
�3�����I75���2�N��B����E�;u�	�b���U��w�q��NF������&�%0�����st�ګ�%`j�L.����߳%m?�|�92��Ӷ�L�g}�Fay���ϥm�g���=S�W����Ҟ��Í96&�Pp{�!�I1��wv����zЊ8A�P�y4�m%g�x��v�=@3�Ɉ�[�A]����&��J�TQ��|���;b%���vd~'��߇i���1�����մ!D��N?��]b�-1�U8��H����r��t���#Xb:y�E^�zp�Q���@�␿'��1���/�Ul�������jMfT4��������Y,\ú�DnԾ��m�x�(�˲�2m��=`�g;2��zx�痪���W	������>�.��f�~k�L��*@#���� BD�n�m��Є.Z���s�ٲ�l��C�"����3��]��vsRIOa�0jp�n7�����Pj͞<��\��e��~�◡{�J�2�I!�I�\l4� /La�X�*]S�f4)�%�Nr��CCX��T�is��&",6���Yc-���Q� L��v���ڹ���p[��F�m:���vK�����1�~���� �BVv&l����*&�9�~1ro���@H�F+P���Ěf0 K�$����l	e����&���MX=�5��W�0�L�W�	5�閝`��N7��I�I�ā��6M��� H}��Si?�,h�1��	J?�C�X|||T��U_��3�\`}�{Ͻ1W��O�`*ۦ�6�Bd��{,MA�Te(�Q�v��w��G�Z��M��Jb�`�a�nM����D=��9�b_�(��}n����cڌ��?e@[0�sIc �y�Ǐ	�~%��؈_�se�w���c,~(!F,�\�n����w{�1M�5X�X���=����yQ�渭º`�'�#�&g%�c��*��o�l��J 4���	@^�Z;h�7pe��9������9NVxJ�6"-p�2BP|��Q��Ć����|�_��p� �k�!`�������yZ�U���F�^��n�7�*`��U�T�F1�z*Rָ�_�u\:B�Ⱥ���/5_Q�V�̆��0�è��d����FRJ���3��3Q��u��$j��'���6HGP����g$�Ǖ\��=g1�Ւ	�ݨ�??x�3�e�_��
$d"`ȯ��_�8xOƟ�k-k`� ��m TclF�48<���c�����:�T|'|F����nY	�8k'1O�M�&-F�eYp�x���;��Q5���$��d��i��۫W����a��z��.���3�ٯ l?S#U����&խϚdp�L�~��$�iŹ�grغ9p=����lھҎS�f8�ɂ�6r�Y�O�yf�I��:�K�C���t_�)T�[4�;_!Gm8�����3Bk�{�4%�1`�����}�ùm��y����*|�yD��V�+��+�=���wp�MN`WHp.-�����!�1�z[C@@V3"�����꘦�S��)� �km���7�tJ��y���j���Q� ��<��
M�)���6�=8V�0+k�le�K��
�/���o�}��-��fC��4��6�(����V�l$�Z�nS)����M��ݽ���sJ\�`YfA:�Nnr�����s"��`_�Rxl��A�L�ٶ�}'��]߀' ���?{7Y�'��yV�R�?��v��{]Ӑ����v��x����Y��K��Qy��;��MӴ�JI�d_�g����f���0���0x���'�?>�������-1��du|��!�pZ�o<�ɐ�`�Sye�����V'���/��ŧ����R]�o��ÂTj<��sٴ��5_�1J�����w�q�"�?�IS��+������=:�mˍ���ob8C�ir�q;i4���=j�^ڳ��Z�o�zz匰�#�k�O~�st�{��zg�<�>r��Cd������h��-�;����ȯ��ϽgYMm�הׁK�xdnhהCe#��Y��\����e{zd=���S�ֹ��O�-�>��%;�c��O�8�i����ۿS�2c�`��& F[� �E�	�yDD�%��7̏dCa2�H]��zB'�an��ɰl��@_OP��T����\�,(d�;�T�13�)<�� X��ۍ���<�/��8b��u��S����H�i�j�Ze$��&?8/xN��w1Vi�(�sn=]��������Y�mO|�ގ�>y��r�M��Ϊ�G�[�P��~/Z��q�}���&o�y�G��!2m�5���Lp��*]�\r�߫�l.ό!���JY�9�q"ͬN�,姱��{���7��-� �J2�E��S��\î��P�D��c�]oD���:Y�5>��5!F73)lIZj����|�H�Tn�w�,3��}R���Q�w$,��=�*���3�`մ2�Wz/4���OsgYB�X!������_��jQ�.3��G Tޫ���\��lYT^�ݟ��j=��3h�i6'�U��g��eB��}���1��kTK����y~uh�g䕇��RsM�w9F��'`����T�&_�!-�����|��O\mb��p��y���,�,�4e�fᬃ����&m��oq�����?��ʳ�Ex�dFLR�͜�jrNU��`l�uD����%�<�y�n���U����v6��n�S�]_��ɚ�� �_�����h���Y�	;Dc)2�Z���#l�f"qF��D�\qn;OZ�H�6m�k��=��(���՛�jR~'?�6�BZ`���Wm}���Fנ#�K�{���-�;��)��dҺ=veh����|����&����!�D�%.0��`bT@�h4ll2�F�ծ���d����ZO���`&c& ZP���s���>nn�� P��l����8& �-����Z#s����C�Z��,����Ő�E��Թ�0�D}`!ڪk������i@W˂SO��\�!'*kuOP��[J���Sn2�KT@����}�Z}���f�Y�W@�����f:�>�.AD5� �,s/��c�zu��_�]��BH�1��g)�^(�T{e�YZ�k}̿kZϊ|����>��l�6��|A�ߪ��f��i�S���iL�mI�@�f�ɽ������^�6�2�h4]�������[�=��J��?�������f�2���DsX�'I�yF�<c�gx�,s���b
#��}ZcX��q����;�kr�*��m�{�os�1� �`,��@�O�g)a�SX��u���Sl1��M��&>*|�������XY��������j�9U�� !���Q����Ł���@E�=ǞnX�w-H�l/��h��d;b�a�{�+_�� yV�0�-pԻ/� �u�(��gt�M#����$ö���g5W��/�n�T;r�hLFS�&z�)�kʡ���ãR�MXA���2�e2{��B{��/`�o�~�W|��~��~�c�|��[څʹ��;̥3���A�&�c�06yn�M�.�"�ϸ��^d������T�y����a�eX�ȣuˁ֛\-&!}f���/�{�H�6<��;� ��b����E���s`A�ʅ`/^&��!���ok𮱒�aiOF�#�:�U��]G��dNt��Z[�����9��&!�&������(2�����+�B����� �\��N[�^�}�͊�գe��mF^_�"���ۿ��iG�0�Mv؆�"��1ʔ�m�A�Z�J��hrM_yެy�
h�R��d��!��!5t[z�B#�C��!ȊE�ٗb*�b�L�ʓ��{uJ�('����Cs�P�f��WI/��j�k�1)+N��v��ț	��뚐S˕�G*��C|��1�WJ�Fj��v��k()�y��KȌ]�m�T��rRQ9?#GgG��~��7جR��a�����I�ݥ�'UxRz��g�q�0��1� �`B2}�h  ���swՠ(!�욉hcN���m����YkqD�^�s�Q��������;�FćP�f�D�K_�����%1ƍ���y������[@�d���<#�e�6�by��^�Lk���c�M�Qkm��} �[�#��P� kj/o^w��bgr�۞Mo�����k��ۡ.��O�y)gD�8�,F�]���X�0	�W�i�83��کL�x?#f	Z�>�d�=ǎJDc��h���rBv������X�l�n$�x��3ND��*$��Ѻ&�چ�y�y���z�>j�ؠ�c]�{e��}�8���%��M�&v0	`���v�c�g,�����i*s��1!F̿~��~+9��5F G@'?`�T��)�g��cz+�e�	9#g����,G��^�S`��
�%���i}X���J�}���6+{���qu~s�Y�%�iF�����]�M 3b2�3|}?��^0�=!�r`�1΅�سa�TG�^)=�h�9���,<_#-���%F_<е�B*�?��BA�"Ν��b���V��>�ĩ��Z �FĨ;��R�FOኀ�ᐢm��@Ӧ���4�{_6TM��E�n�����F�Ի=S�_�~6d�\����f��f>A��ce�Yg45��`��X*W�y��.0�<P�f$�Ŗ��٬II�Q���M�`y�$&���,JL�dO�☭�+D�F|�y��dF���d�e�ןmƶ�(o���3��?�'n6�cr�1$�r�\D�CI6�c`���D����	�*ל2�L�a��`���4l�櫤R�F�'�Z`Uʕ�F��
`�td,ˈj�l�VYb�>���0y{u���D`l�~��.�c�G̃��V�(��J���9��Q��2۫����#��c ����l ̑1\��	HL��sjg�y��gu��t��C���Z����=�2�>�J����- �O�����?��X~�	&θ��/���� ;9�yƏ�@���%���̄�+Gڻ�"g{� ���=��C���M���V�*�.'���Z�%KPB$ �-	1d6A�3���;�>&q̹D�)� ���496�t�2��[��d��J�j[K5�<�^�{׼D�c��kOc!�}G�sD~�Li*�3q©��'��i�fݯW�1�s��߃�����̣�v��g1��^��M쨂3�"���PY{{ő�K���h}�=��W�1�m|��X�����- ����O����#����!�����h���*�lN���?�1����� ���O-qA��؛�4Y���3S:�����13��ɤ��6������p�Y���u5��Nr=����R��L��Eeo��A黜vч���b|�,�@��=�����?�"O�2暖q�A���{�	�>�2�bV�������Gg �3�XX���Fo�����7{`N>��];�6���fuh�2n�T���2zϣ���gF��F����N2)��{ui� ����lj��:���%ߍ5��8�e�i�^]"m�{�H-��~�s(���Vv��N�}�W:�����y���"q@8­l�4ߚ��4�9�e	����g�G�6M����1�����-?1��߆4����^L��B��<򻑷�L3��L~���ۧ\)ts�&Os
uS A��uʒ*m�EŒc�q��	�r�{�Rc�m)�]}��&��P}��g�d0{`��+��~p��\��90HP4Z�#7s�a-[���-A�	���,���1U�M�y`�) �Y���GX�;"=�i��;��w�T����bL��бSG�X��S6h��o�#��F�_�P�3��8	C������<��1�H���
�����P�h�zL?�{��&3���\o=�a�ak[����Vl�2������/0�,l��.�֤�R�hU�Y��B���d�:����a�<��"�����6H�5\�~^��o�\4���@(7��3���RV�����8��B��z�h�g��@X�|o���YdGU���{��k|C�e�w�<�,��@�2�ƣ��}>[lo����~�%��7�ʸ:�E��އgăd[��^8CY�O�#&m ���ɣe�0<������gm0G�M{c��u�>t[���������.������{��ϟ�~A���O0�2��U��|"����xꗫ	-ĴO�}���h������Ų,�n��{�p���p��NY��ݩq�s�JY&�n��,��cY1R;<�͛3��"G�ߏJ�	"o]j;RNii�.�ɘ@�:�1p{�����X��4������bJM�7�3l7�uk�����ۨh���k{�ۮ^�G�'_�y��Qon�nͤ�����/�F0���mJ��uί�Gg���=�"�q5�=�½��eAm��ެB��vqGR������`�i"��ºB4����A�H���-�5�H�"Zt.��,W���i�mw Z�' eq槽=BX�Yk^�-��v�=��P��ڪ����Fn<v[�GiLu���m������%��%�3N\���m��1I���4�J�q�H;1�	� fjb	{R�g�I�o�e��ٹg���&�ZD%Y�U���#�~)��rk�}�lmfs��ȁ[c�G�:��V}.�-Y>|���E7�i��vm��#_7������U3��=�̡��L�w��� Α�$�t��8�k�6n�T��
�ɮ4�n�eb'�e��R�5M�\ccXx!�"����H�k����كVA�/*��ׇ�;*o�1F��D����2�s)n�s��0�dsA? ۄ(;3�����z����M'��Nj�r�L���g�a'�HӾ�ـ�v$�mL��H��1��j!�7g=ǯ�g�c���tZ�э���Ku>��~�^֔�\���=G&��߯��޳��)�F#2�Z埽W��&W��-��;���Wm��~���מ��6rX�U�ޖ#�M���uc���~���aӏ�8��E}v?{�~���^!�Q��8M��L7w��@�ܣ&�F����`3^��m�n��5@L�H��{l-iyas��r��f�ФB�
-�*�o�2g�M+�Ơ�GӉ��h~��- �&e����z�V^�{�V�������+Gʤwƃ�����?GXޖ�g�sW��O׶�y�m�~�^�Z�j�x[�h��C-�`�2��\G�Mh�ߩ쿑�����C��q�&q�;�rO��4"�U`�}w&�Yyȴ>�!���8��2��^R��8��,�቎;ճ�l��.k]Qg��K�p��A6��/t��-s���!�B��OWJ� ����L�	0y�c`�[\^�Z���6���SB��,p-�#*(٦��B�l����s��D�ά��Z���h_�����w/��^���������~�|�wT�٫[������xf��9���1!Md�Tف��q�ؐkقʺ�c���1򈌂���3�=�8T��ȁ��1C�����gذo(o�w���nr�m�)`1��&�5l��ʂnL̋�10��Ā��dX�x��mi` �,�l���  �s~`�"b����䁉k[�=�}_T��b�W�m�����o�����E���<b�wx����4�$����D��4��i��,-�F--�?�ܴ��46�V{Z*,^��:��r�4Z*WR��� e��Ӯ�ek� 1�@ݼ�Ӣ��d�y�h�����;�c��=<�g���^}#�L�0^�5v������L�]cI[��`ܙ���p˽X��<j[!��1@���Ȓ$tj��[���6j�zm�hi\�xhA�u#�w�ٌ1)W}��0�kl|�X 8XDxX�L�6L�0�b2,\�qp@�	���c�6�m�C�+�S��71�S0@�A_��D���|o�v�B�z�ez�9��A�=���#s5�ٲ�����7��>�[�����A��S-1�~�,�e��v�!C���r��ş�5��lǎH0�-�����[[�+����M�U�\3F̞P�m����N��u�H�sT�CD���{{%C���[G�%GιQ�}T$�Z>�i$��J�~o�]�4��:C�h�9H5?��M>W�ۈ��<:\*��Ɩ��5��/I��]�J����ԽG�
�+B��f��4{���m]���F���B��rM�V}ZB
i*�g�l��`�"r������z$C^��>�$�'���1�Ē P٢8j����=G&�������]���j�m:�>�1ã���x�zG���X&-�ճ�!1}{lf��l_���Yq��β&.ə�/EzkP�
UEc��#9�&i5��8�K��[�����Qꬉ����H_<��72]�B��]��i��	�ž���!T����]K�tV�į�������R]��H�헱ئ�h�n��1јŞc����E���s�"����͜�.{�rF4&h����2�@�4g��j��V�r�xn�v���hKF�ј�=0/�&�D{rt�!!��h���m�v��3/�7V�hcs�^��nf�qu[Zu�l�Fu��z��TR�9k�G��g�����'zY�F�bR��_��_���dr�wAR��Z�Y�fr�%����'�1��5�v�.�_�i�8� ��k ��	�Y�28B�Q4q|�~�ojr���+6��)0Mz7M�a���ژ�C$<�o�p^�~��̂j�<����0�**��Z�%�R�{��&h�fC���Φ��H\4�٫o�&��e�]�� �S���OT��{���ی2r��̢U�F�_m��T�{sM�K�|j�M}H�K֐�9�z���r�q��:T�2z���>Z�����u{t�n��eb& ����fEcf�5I�����9���?K��;�vgE�f-k�'`{M���_��i+ư&�h�PS�3S�o-���LS�w(W9gI�e�k������l���ۘL7M)V��`�;�����i��d�	��X��}yi���{fRU)��@'��S�~-�qX�Evuq]��򷶝֘��#��+0��^�d8�Qk��T�������'l	M*�y�~	4��)�X�gEۈc�n
�P%X��0��/�i�)]+Y(	
_-�m���-R�bt_-����a`DZ��+E���1�e�V�go5F�b�ͱ�W�:W�A�|� 7�@qk�;�\-�>������k�I"(P�zp���$�:��[�	[_!�����_�������B��)P˒�LWk`�A$�����5M�QM��j�F��t>�!�F{fq~&��hk�&S|Y�ȎJ������-���F6�h�l9�xjR���
�x(!�~�<�*�@�����r�&9��1/Y�=�q��u�ɬ��ki����~��o�H���v=�~�{�Z<�f��^[\c|���}���w͝w4�u�P�9����l��X�#"��U��M����8Rjgm_4�az����֬�f�ڴ�|����C�Stj1F,��<�d�2{�9,���R�xXL :!n���x<��P6w�,�w�ba��o����WK_U��.hm�
��QimΪ'b'��,_T�<�����@F�p����Ǜ�O�8�&<�On��b�F�������%������&�?'��8x�ͯ籭�A�<%�eR�`��-���1����^^��ث_�Q6�+J9n���-P�����v��=ϼ֪[������Q@�'�x�#f6Ƭ��y-}ŴR��|&�Yi��ȡQ{'�^m�@��Y�c{s֭���[�b
9TB5�
�e��}Jg���L�"!D|>>q��K��=�/��f�nT�v���L4���z>FL���3�g�D����L@4S�c��X}&�M�~޶PN���3��f���Y��j����$L��1�	��0�a+�-�bۘ���?-�l�Lѧr{q�8I"���_�[���TjcT/�֦����ρ����P�l+�2y;F�#A3�]��N%=&Ok������nXRZ@v����vK0�����{%��+��Ed{e�����>�`p���e�Y����$/ս�yժs��%��$�*�XZ�r�%z(k
{&�~��(��4�m�g�o �i��H�#s����q�������CBԿ�n�s>>>��O�2Ϙ���~�d�!bY���;ܧܦ;�������?p��=n7�G3�`B4����x�{��	��.�W�[@�	(���ǆ21�De�+�vF4�|K�@m�?s�sd�|V$������˛kL0�1 օ�8�0�#9z��آz�>��mL�v,J��&ز���7�����6������v�6��*���;9:o�3^���AF�[{��akЦm�ʺ�{��J��̀�G��p )���Qo{��H�7����E�!Hi7?(s����q���h�@�=�*�{3O>r�����W���ȕ�L~�:���n�)�8%��w��8��1�Q��٠�@�TôNɚ|����P�\���%��|QCE[�K��#R�MS����,{���t��e_%G�����d�5W�(���${��+�7(�]�T�Yn/��^����K��odm=�>F�-5��2C"��d5G��xb��9{7���e�U�ɋ�%�K��t�1���]�5��%�u�\����W���Z��]n`�M���� �/(Gـ�g#6��L�IB�=����W6)���ɑ�B�p.�N5�U�;:����r�D����6�q���2W:� R.aY��#bQ��g�q�#�·�m�ϖG�b�Z ���ppFzl!�l-�Y枩�����`K��������ޟ�����Z�ѭ6ҳ�N�2y�1�8R,�=��T���m4c�j7��,�w��c`cD0ac ��L�#�RZ�e��˒~��Y�JB䌼�&sY�c��vfb����)��A,F�=�IU�b3A�y�M��,L9� M���Ox������hx4���>�q���E]z�or��A��y�[�?�Pŗ�����a�K}I�,�?~�H�ϭn��[ e u��X1��hǳ�Բ�5>7�l (}�m�<~��fO�q�ϖ�P����Wϙ�[e���L���U^uXuk��gګ��+���ϊ6.��Zij�ց�:�7y��{�E^O)gp�V�y����My��R���#� �E)���K�\�}5!�0Xյ�c�{����f�+�s�$��۾cR]�	!��5��)?w��7��o��	1�3kM���&����n�#J|���;�- sY<�m���`�bڸ�ޯ'1���IĜ�L�����9�/�TV�0���|Y���=��.j0�z@�ݺc(�W@Ȭ��yYV�������m�+�J�y�	�h �6M�t������j=[b��ƎT�ޫ������4 �܅�����}����qL���$�.�Rʹ�9)u����8˶I`Ʌg=*�5ٔ=$h6��sH0�R�����I*���Dj��Vjt1��ID����)���T�m2?>>m���x�c�ĸ,�S@��ں��sf���+6�����.�kH���Ì^O��{�Wf�A����M����v3ƈ�{ܦ>( ���N ��V4c��{}�PU�ُn8U��R���-*X�I&Se�U#u�7�h$�G+�ra&�����v��k�C�-��� D�R�6���,S8
�[ k�Ik}�ngT$ o1�o����m,%����L׌���=��aCk�������H�f�)Yb�:tE���YjMZI�����u�[H�ފ���u�|F/���R{BJ�=�OYG��C���;;m�/N�`Y|J,?�@#�)�`D���V��F�:�b^9���#O���@���As?�MO(� `X>��ٛ0��J]|��l�0h��q�D˃��M���2�Xc`��6�^ _^�N$�h=�[�ji��V{$��Le�r̗�_@���(����YU��� >~]����&���[��>�o׻=����F�����sd]�!�N̦0�Gd�3?��<���Qi�1�y�8I(6�ZV��}/���]#<,�7��g$��db�d`�N��G�s>f�M��5N�F�����]�,��?��  ��=� � )A�`����t-]o<#��F�~7 �b0��I-��=\�cā��s����1ݰ|z�`0M�qi�ؔM(ڀ�T�I5��c��>��cEr��y��o���|oa�'�:�R,�6<��}c;(���U(����veC/u�t�i-ڼO�FO`R��R�8�<����ڀ�gk�����~��e�yt�����.�{ �w�B%�� c�ͭy��%^g���R΀��L�l�&��V*F�V�?{m�I���7t�9d{[}�;�q0%���К�����Ş#�Q��n;�c.��i�HjZZ����� 
�G�@��v��s��<{�Ҙg�w��X@gm��cS�hc�`�Xd6�V�� ���X��4���"�O�0&�� x����/<ĸ��AW��d&�w��S�2�v���@V=�0I��1�h~:O��v��}&2�'��1{d�>2Y[ϻ.N��WV�u��|#����X����@��b\3�H����GD.��G�n��g�T'��/	��Ro3�@��=�~Dz�^��!W�_�P��F�	P)�O��~𵞣U�e ssm��y�T�����7�ߍ�jv�]T��վ9�3�ష�$3҇��݁:�O��+��$φ�{��wv�޳�ާ<����:�mn��M��+8'P[.�3tv��`Ik��`�N��(�X�W_��mO϶z��)����� �>c��׸z���XU@%#���9�@�T��˙��.|���=c�I���7�R��{�HP��J��=�ɨYka�-�4��	�t��:�y�o�������:`a�F�к~�V�"����TC�)o)�z�[�K9���M�~�� �ʉ1����$��V�`�����s[���=��!Zcw�zb��ގ�����p�ڹ'����!���[@�<Ϙ�9��B�|�M����d����joӠ�bTU��) ���j���N�ΡVq��=!f��6��Y��= �߅��kW2d�m!�Xˣ20GT�g�LE��{F^�&K���#�9�h�w�y�l��^��;\](�Qf+���O2SKHS�4�i�ʯ�0���#r��]oi��Lnv�,��j�U={��M��9,�/XH��� �-�����0M!Ƥ>p��,p���A�\����z��`1�w�0�1��Ɇ�ּV��l�1J%��dp[����-��E���I.d�ibZC�`MR�[�2��n`���wƤ8�!$T�F�o�NS�^>w�w'��H�t	0ٳ��[52m����GNYFKE��FR��c<�-��훴�[jޑMO��tx�mo���b�δ�;fy��{�h�-净E�G������v��ɞ�^�{׏ʳL�H{��zg���b���o�Ny�|�[ɃsK�)W�R�+(i^UY��>9zp���W�(W3��a,4�2g��[2�D݇�y�c��v��1����4³��� �-9�~�J�k6q{�&˒��<b�g��`"p"����4N���܊=��1��Qa5Y�~A	�y. s�I�	`o��Rrwk�i��BXnr�p�	!9�Ђ�6�����$�ɴ���֚20Z ��x X�u��j���E[�h� ,��@^r�0�F���E�+֘M��y�gW1QW3Z#a��ZZ`lO6���E,���)��r�3��BUNվ�&����50������׀�^9�v�Ԁ��3��mtn�|��  6��]�7���Ѹ���e�y`u�f*K9t�����"٣oݳE�����J��n�)��=����Y�%�x�/��0!es��ֺ2��P����2�����d�e�gƱ��˜lZ}k�;�%�B��v����3��!9r2K�ieMYɽ�k�3��"턞���Mh!ԛA��C>x�d �6�Q��b���β�/{��_�|e��m��V�=��U�zE��?4�q����'�v�zx�2{�=2�i���܎��y�Ȗ8��[5f=�����17]*�|�D��M|`g��[���ʤ$WiyFD3�1J���Lg�8�1f���}0iC��'�b��x���(os�	dlj'�����F�!�`���Mo�Uձd����;7�	F_������d���W�/G�T"-���'�>��N\=���9��4�r��y˾G�e����Re~�=��Uh_-�m�\){��}We����Zm��y5���C[Wz���+��=��y��m�-��,��U��Brx�{��`]�Yz6e�%�C���⛸��n�aP� *���`��=c,��-E��Z�ƝAk���e�j��ٹ���gߏy��9?�+����0�+����Z��s�}^�b�ub�7�|����p�>`�����'���`�&��5X#=X�R�K�X�9�%�E0),D�44Yb
�nV�6�Dw�	7?���^�2ψ9�G4��ƒ��'�FU�\<9s�f�jU:e|h�zh�����y�j�l�q[����]�g@�Z�����Bȃ
��jӁb�D=f���f�R��6еHij]y����1YG�y)��Z	j
��8{W��K~P�ګ�W�v_!G֏Qs�#u�LQ��Uk�r��Z���*u\��- w���-ױ��ߒr���i�0�����z;�ř��(�fOB��??a��H�T��<_i7�H5�0��Me@���kC�X��yɦl���uN�>�����B8p����v�����v��_o�]#�9Z�:��w̟ܦ�Ii�����7k`aq�M���X��O��{�{  ,�^S�k��S��������#�k� V0a���Y��1�l�<���)��`�xp�-y�%��l��&�+廳O\%��3��&�V��:c�j$O��2�UY���Q���BQy8�h# �n|w�ë��*`J��jm��m��k�G�?�4&���]�K�8���sn�~�ա���������rq'A��5��Z?��H��� M1�z˞òn[_[�
 J@����� C���m�g}���M*/��c/%��޳S��'�k	?Lm���r�'��Ȭ�5�&X�fƒ�$	oؼ���C�d)���)+3�K� �K�c����7U�D�h��T6z�V{]حs��崒��+Z}��;���$��A�/9�;���-�9�I� ����F�A4��4�/��4��V���+X�V�Z�����B s���ɩ]���Y�L+���@�Ȼ���JƶW7������w9�2�-MBk�HFp��*G=io�r��gd<�;�4`kYh�3 �̭dE����Lj�r�=��K��9�sz�F9�E�q�!"E�������ް)�yظ��c7�����G˱0߄���d��i1n�L���^Эu�ԑN�<×(���geo�&��&��f:*��3�˧�bw��s���^[�m�;'uШP�P͈~d���<�a˾L�ОZO�uς!Y��8����[ԑ�δCج!$g��� [��u�^�[��q��ڿR8s)��+̇dy�F|����"���CR��\K����V��x�uw�<�.u���g=t�gkX~���kO�g<�Gi�߽������P�p_�t�B
!�=����DD�tn�}��8�J ����.�`�K���ή�?/1�X�l$�ᶛ#�^ �*Tʈ��ޠ�e�끊���RͰ\����	���x[ʿ,YB���;�@�)���yD�Ev�1�,F��0/��G{'f�Y�PM80���yy��Ò}z��:z��������'եϴ�T[ ���1�B���c��;:�{��^[��}�m9R&P��;�7�ZB �k\�����p���x<J(;�o�Z]GU�R�9�LY�8�@�<���^�٪���ᩄy�m"��fo9M7�V�1"#�Cw���X�އ��Ɣ`�-�<�#��ZR�Iג�ni�X���Ѱx,~�����3� �f�Q�T���5NfYd^�	@�%{��>n���6R���ǔ��:����Ѷ�m\G��3"�E/$����.4=��T���;���H��g�B֋b���|�;��0=gA^�I}ٸ���'뤨-Q��L�߷� ��� m݆�ln�� H^b�� ,�Y��h�02
G�)��gAߞ\9~�?-�hc5���G�����
¶�i��Qab��z�_�'W�Y9����[��N^.�&�b�&t�A�>9�F9o�FZ?��'�3eܧ��uZ����dJy<���&L�T�GŴ��Β��L�b1��֧��@C�jR9ɹ*J��[� �*�q��ը<��tz5�6��2�����'�H��A�Wj�������a*-�yY��:������F�6n��2`�5T.]3������8�Z�G����)쎎���G�����@�0�$\��3{�\�G�v��n޳}��d���ɒ�Jζ﬌�uԤ9ǭ��f�T�9:��&;u�I�o-�8�<�<ܓĸM{�K�,��wJ6 �2����m���]&��En�!}@l����[���C6�Ȑ�ɲ���/K�˹������0+��Ar�yq]�4n�#�C���������2M���{g�o�>y��]����ҋ����U�A�s)�\�6�M.� S����q�j�j� ��@��bR��}��ZR�+�Z�H���z�~c٪��������̤@��:F�#��9W����������gr\�;z(�}���;mjC�^�8�&U�F<#��t�x��v��r���V�Ϩ��u�~�J�Q��T֞Vnt.��5�~�)��`3��[r_��cH�p�Ӕ̦�ɜ6�RR�M�}�d��)�K4�0�ٸ��fHc���2�Gy���7��C:������I� �,�8�3ƈ��z����"c�0�)���: "&����Y��b��1���r�������~*��e��븙�~W|[�g}һ�*�⳱�����Tw�E��in�$uDf�3�lC�6�����ze�T����q���}t=}��0�KrDrp���ǤL�'�xp�Y�~y���(�1��^�Ӹ���fScO�6J`2
�G�8y��:�P���ƵF��G5N����1!s�P�o�pH�z�Z�z��&@��l	�'�1���i���|~~�k��.�󢩣��3�b��Y$�I�v�5"Ԓ��ֱY*��A�Ɖ��Qhc,~���Y��s������2l��!�Ǐ	X��b҇D��ɕ�4t)1�d,LfJ�s�&7a^f̏G���3L0���&�qw����#��|�ۘLJ���j!Z@��4��e�<�)��<�v���!�0�źѳ8kV��^��N�Z�ʟi����Z�G}�F����bOx�`Q1�<��t�-%�f��}�Y��������v �S�V�TdH%	Tz�!scm�P�hϫ䨺��~�2/�P�qtPl;�L�� �fSc�5�,ǀ��(��ߟ	��:0���+D�?Yw��P�=km9��v�CX��������Qƛv��Ɠ�!e]� y;���Ѱq��C
����׽�l�a�g�G�`B��6������-!{]�<l�H��:�{�YL�+j�a���b��a����~��������������2�9��'�&��X�Z�o�YC��f��O6�����TN�l��<�:y���yǵ:{,�FU�m��+��U�����#c@�l����mҭ2�f�﵂��{���w�.1F�F*��8��T���Xye�\��[��=�s��{���9^v�ܫ�l�B<���@�]�.7�H�f=$H�&�F-l�~j�#cR;<�$!)�I�i����"�wY��G��X�V�h����y^*p�L���n�0��7� �kq�Yy�����o���w�&�n78�p��6�[q��g��ނ�euz�3a5�<-�����T�s���8*�� ds�N���2��Q�N�2	�_K�ƅ?KO${�L`U�I��M ��r���l��{_������때c���.ǈ�8�p�WV�Y����u�h
4�����b�|�ki*4�3k�ޕ!Zs�S��Ϭˣ@�"�[>���\�@M���k�3r��g����j�~}���i�0x���Q���GMFd;f}��q�̘�hT��d��-��b�|B�.��� w;,q���'���}�������������I11���,��]�/>���y����ь�����IjZڠ��m�r��"E��� �p~�ֶ��Ƣ!Ӧq�Q�@�1�6����v�ޏ�x��ɈzS�?�5앯-��ѭl�B,�B��˲�rd[�)���{�^��ތ5���� K�3��큊� �w*�q��x֓;�j�Y��U/S>�+�m��ֺ��h�7�����ڵ|��������F�<-g��>9�{�v��R�*��,�D�9l��PH�-��|���,~r~e�#҃����Z76�_\͵n��&�ё�la�c�}�F�.�t��&�#Dx�1�3L��c���_�~/s�����\��9̈q��Fy&����$�&���.��B � ��&�i�Q�Q�fc����э!x�(@�5f��b�C\\%|ѿM��S&��8����R���b�ɸ��1pVXu��N�����fd�	`��SμoM��w��8a:�1���Y���M�c���u����!�u��������C�ݴ1Vq@{���e���$5S)��>ց��f�ٙS�k�\�1QkPlS��G��oYP=W��>2��¬˲���r����e�����#����ԯ��]�̖:�r�oDxư;�Yb>:�Bx� ��IlP
�:a�Ȗ��i�(z��N��r�-�WMF��H�C't_\���k�qM�X����?#<X?�����6�6ӄJ9�Nծ=������w8w�"� ��|��V�$'�P._��:�����
9�^�G�UkVa-J@tn6��0�F��rO���VcV3�M$n�u����G�w��Y�$0z�n��}��X�� %�����e��#bA�b�0��L?.m�3����]�����~~���ѩ�7QL�n�;�eY`�ò̅�;㹹'��[
�L.<�e�A��4�*�|���V�q������L�M�!�uS,S��@�F�wl7@�Ik,�(It����</���זJ�'��%�@�9#��^��z���I�g<*�6��%k�� ��{%��H9���Z�Ϥ������K3ay�3�!�ʦ�,��E�I�vR]���z�y)�2� mrҌV�ku����G��6K a�|s��Si�T��� ���Z��bk������t��ly+��v�A�L�Y�n~� �5�"Vr���*(���{L��'�>�� �2=>�o1DkAF�l�����hc2c�0@	�`���qO�z_�(���`Y|~~�E/x��n��,P�ӤzZ�m���[3v|���2hz;L���٦�H)����H���ևR���c~���i�U6���#J�p���eã��vq/s��*���t��Z���l�?�4aY||�ՠ��*�����D��r�"��e�2fO�;�>M���������4k��p��U�"���e�PR��H����êι
d��9�[ ��w���޿��.���}ڽ1&p$�;����8��;�>i?����Ekg�{.Zb-;�3���^�5�+�ޘ�����2E0����KA��QaKC,�րD�H�+Z~΅,�>z&M�|�,D$�<,X;��Hj���˼��>j74�n�����;�	�{s���o�1x����#vsƲ<�7,����w�;��	����Y�����������L�����13w6��K�~UE�K/j�|�X���5��SX���������ƤX[�w���Z�ۚRnmO�tgCo�{6Gpeq/��|O�J �k�T9�{�j�r��r:���lj��φ�#l�(��׸�֓>�@Шh��+X��pV�׭e�y%�ə]u������|��@#='�*�c����e���*�non�MC@�(6��Z����=`�iZ^%�&=*B�j��Y#,4a�G���^b�cX�@�=��D�O�<�id�
�#�s�v�K���X��9�p�Mnӄ�M�n�J�IV771��xտ%Ud��q)6�����~|��>���q���忄?����_�_�����_�����>|��)N�3���te���=�1)�d4��D~i.�r�I����K����q�6 ���ee;(�v���ϸ+��uYĸm�4�n-N�[�L�S�\�\������Mr�,�=��a�IZ����e/ړ=�"?�n�& �j��ٺ^�Ei�H��pRUzD�1��e��0F��QIj�v�����{�ϼ�ֆ\��������GD>+��{�s��(o�wb0�����,i�b��]�N٦}<���ұT/4)��WH!�b���&C��ަ��~Y0/3�e�<?0/3`��������������������ݿ�?��t�w�d�5����&)�`�TV�ZL.�ļM���&W��ƶ�}��D�oUc{���ސ�j_)�η�b�1�P*�9|��ϙ۟��	m,�%�E�!����we����GqM}�R�V�̎=S�ٔ��~�)�aF�e��^�&��}G��
��C(̗��^%-S��q���a�d�m�/Ǽ��(c���������)&d$���CBZ-mܵ攦͸R�1S�R2�l��g�.m5�������iY�1gƹ6Z�P{��#��Sh���i�*s
�H���?/X��e^���R��n�oR+[������=���0��e������g���<��w��������7��������_^�og�m ��}����f�x�W�S�&�K/�˃�-TIn�in�;��;n��/_8�e�j^���lFB澵Xf\�*��S�l�n�,�8duv�,2�驘&��qġ�ޱs�W4���6>�����V�H�B�oiW*٦S�ə��H�_��j���o���ɹ"� A^w����8�=����MV\��L����7�Lq�:���v��#��9/ǊCT���4��4P�z�ʱ#�K�g�����/��R�[�u�n����u��G��s�i�K:V��ߘU�5��J�4h�<�`��#�$�I`3�[�q)LY�x��"���\ ؁��.b*���������`��:��1�&��o������vÿ�����_�7����u��=y��j�-�%�!�|��K; �-'O�3��\ܾ����jJ@��+�,n�H����t�֧���e���Q0G�ܳ�BFA鑲�f�����
��a̞�o}��W��+���x�{Ř�e�h	���^VZs~��u�q��#m�\��J��l�1D,�G��i��7�'|�o��ɤ �Ӕ ���XI-��49�2+�c�f܍��Ŕ���<>����gLH������d~������W&S�Q�_�BFOH�'��/�����r$C�ڢ\	�Kؠ��(�=��K��n�_�5N�C�c��:iS$Y�͆�Cl�y��J�ٻ��pM�6Ҷ8<2�2qgE�d�J`�U`��It@.G���x>[ޕ"��������j�5l�޺ ���1�l?b�|�pu8�ϵ^Z"�w2�\
V��V�Hf�L�I��`���`Ln���ƭ��1Ɣ*2�#��� ��`C5cfR}�Y|1�C�`����t�?��?�o��^�]O˛���w"�u�L<&�b�^J�T1cy���E9z(RSQ(����0��"��l@�-��H��v�f����B�St�%Kgiqv�0]�����6�d;�wtS�0au�r��L�����r����Wk�$��!������>4��!oĄ�'��W��4w�枴���7�W�u��T�Sx<��;���j�e���]!Ƭ�Z"m2�GEF��ea6R������Đ�� �n�>�tdB�	�{���B��7`�a�CdX���������7�]�%����XKF��O6�����#�ʌ��� .�9$�ia��N��o��+�/6��ǯOܧ�%��* `	Kf�r���
��T=�r��x�ɴ&�i�H<�<|���ʢ"`��@	�����̯�����|�ݖhU��P�ݓ:GE2)���*��z[6F--��M2�Rٍ!�n:�z�_h����؟)�H�I����z�h#�P9�|:S�n����������S{���9�Κ=��%�^��{	04`)�E-�{�JЪ�]i�l�9��&-������k�S"I�#"l��i�D�uy���b�9nB�CR�?~��5��O��˷p��6����B����y�I=�l=K)^&"��@p���b���xd���9 U�[� �h�1�(��mL&����F �������,���Z<Z�`(Y��U�������٫}�q��g@!ϽOv!-�f	����C���PYȍA~N�����g-y'#����g6���*��
���JW0_G�����N俽��|}�� 9'ϔ?
�eb����Ɂ�t��W���c��Vڋ��[q=��*�"� {LR�G���θ�����3B���D� D���aY�y�����K&�"bB�00���?�������㋺ⰼ�&���l�
�)��Sd
@�Ʀ"5���dp��}^)�\��v=#����TL���K˶�XS�yR�7۠0���NK��������Ŭ����2s�������P��'���п=���&{��;��Z;��>�z���E�e;��(�Y��v��2���.�T����v���[m��I\�k[:kҺ�ﯔ���_3MS"Vb
�.[�l4Sm�,f��U�~BҞF�"21�3&��Ç<��D|||���O���Ƿ1��\S��)b�R<H�&Xk2x�>�v���,4o_OE}��3 ]�|�҄�6�����y���U�m�3�.��x6	`����"�_��Ǐ49s���mM
�oF�@����Gh�H)�v�K�椓a���۳2z{���
=�����w����rlo揵)$����G��3����mݳB������Iյ���R���z�շ�^��(e�n;s�I#b^�㰦h6�6�L�f�Z��C
�8�.��'e���3���a���G���Ox̳�X5���n���C ����D�* ȴ���ۧ�ҺyL�SRAnի@� ?��~�-/$ibߦ[a�䢛~��Q��T��8��״ �ى�bRC��9�׳Z��	��2��&�s�����!��.���P�S=����W���V�{6m J��3L�f �������P ���<C�G���2���U���ji�h�K��b*_%�P���|��r���6�)te���؊����h�o��:����'��<�"˓�0��/��m���ڒ�)i.e>t�*߹:�V��:�d�:�fY?';H��m�0�>Ԯir��(N�6E��������ӄ`'X�7k0����cm��������^]���;"F}I����S�VL
~C����(�ڜ� � ��s�1eb�A�<� d����p��E�3�l \�e�s���w,���8��Ŧ�k�$��n�u[�#�U��P	H���廳\�`���GD29����c (�m����1s�ɼ
��CF��U�5�$��"^�|_�����9�̬�f� ᶎWϱ�I���=mP�i%!0Ĩ&�^�@���fV'��pR�S�P�h��+����1��P�C3F�� � ,XB��1�g ���q3����%�4X�e���y���R���Q����Ӈ �XC�� {��6{؜�9[�7�1"��Y;*�_Hq5+�nE ?�'qf�6�P/dE�T謅G���b��C
H<"rѦ�y@��J�S@A��p���b��Z��$,���9��9`�7_ٟ϶�H91ƒ,�H����w?SK#0����h��+D���yH$�>xyƘJ[����?�{�*jN���(�G��|('������F�$�ve�H����F����x z*�*I�̞��Vb�ů�w[�5wy,����� �Hr1�_� ���XXc��?�(������q�^(o�.O�`g��h��E#�x��8]Q[�
B2���1�L)����t����讀��Ŵ,Py ��R����|��L���n���'�aN�E����$w8�RL����gnB}t@�Q��zO-&[�s%88�zm�7�k�:��{h�]��m�Y ��&���S�=Ӷ#��:�A�����rF��޼Ү�w��|����0������ȸl��Kk�oXr*��2��O˦��	�`���P�`N��_ß[�������l>��^�����6���Y�I&���;ڔUƐ��V�L�pO@�d�wD}欅�\��\������9��/��y�/�e����1e1�N������'�	���h-�MN=6�M�����1�>��-����w�!�TW�tR��:o�>�c���~��bvZ�~W����E��eh����eAT�n�Iu�ɬMzb=�O��׏��K^v�6*%m�+p/�jiccӑj�^����6cLY��H5�/^ؔ�}�'���Xê/�Oh2�TL���i*�T|6Rg�� �Ֆ=�s��ڻ7��5# �:|�؊�n�<���Ǽ��6i�A+��k���*,��8�	��z�^�[�Bk�<�i77���:�;�~~~V �_�o���3�u͒�ˡ����J"�&5~+׊SJ%�{�<�<d^?_` ��=�gK[�>���Ƥv�&���g�/b�,'�h� ��L7�%�N7����1yy?f ����Tl�*ot�~�e�#\09#��İ`���	�q��4���N���c��?����ng~��5N��4�%���P0��O=!X,~�L\��j���5�)/�)����it�B;rb�>�6/;6&��rr�����&�cǭ�bDx?���Z��j�t��Sg��hK��������M�=¶�6��F%�+��z`s]!����Ū��϶�U,�W0���[�L��Y�e���Q�k�����^�G׋�k�'������p�ɽ�55�H}�/ ��=�JB���W���uǓ��#���s�����:Y�����L;�H�%�G}�'�}B�d�����:ش��1?9�`
;Dl$'1���)���H����L��!�ä��y$R|��987a�M��������/��x�+��j�� ���T�)��:�׸�1ƒt�<S��vzf�g��6Z�8�Q�]�������e��b�N�ܫVc# �I6B`�E���goQ��_��i嵘�^y��J�ŗE��a���� ms�;����H��ݞ��؝�]�>C�1�g�p����5�:kbz���:Ƥ�$Ƹaڏ�ƞW��u�����a`e���$�A����d���rܖ��9r����)?��H�;�;	 V,/�ҙ��y>$u8�=$�B���<�eN ����p1�hC�c\�)l���/�����&����O�]a6�������;��}Lf|Hn��HR�oUz�ZX������s.�1 �)N�.b�n�V�^��_���d
�Vy�c1��`�
a�xTOF'T8�/+��`�s��,��b�l��G�N^Gc��%��.�gճ�~��6WeS�6�+��J�'�߼Zun����?/�T�G���3ԛY�OΕ����GD�4�!�Ò>��!Gz��2�xN^֫h�q�h�������������z�1ZF�٣=�1M��~cļ,������\8���l�ʩ}�e���Pg
V'1c��$���(ɿ��������^`����AD�dc�0�v�v��]�1�s����?��W����y�>0Mn�0M����Dgs}6�MR�[�Ik�]��&L�n��)�˙P�=�ɁbSc0�	�M��6F��1I��aO�y��|:+v&��!�6-�T�F2;����!_�������^��;���Y��yL���[�����)�g�bS��t
���N%�� �W�
\H�"aڻ_>�+��|n@U��~<�_�xyڵВ@�gn�I��A�9z k����z���^������^��kG�������]���#sY^�BI6!��~o$�� f�Id��������0�X�1i�\@�u���S���2��u<d��M�H>	��O,1i����񱾳�ϥB�H����_�݄������@�O����`&5MBa��~L���;�4 W����(N<�%���@�ja���Zn:q$�!���:�d��Nlj�ZG�b9�6�9�\���F� Q�<t�4�I���I�X�5#��lׁ��F��d�I����&��s��p�I�HY)8�
 �烒�pl3 pv.V�a���=�(^��m�5SAK�$��y��V�L���۳�yY��3ɒ�:�}�G����R�W3�=i����ҫ��]hh�*u��OH4s~$Ff��2%�ْ�m������d2C@@N�������,v1H�r"�|f/��e�.a����Iޔ��g[�d����T-�#�Vo�`a��j�j�`��r�s�L)��\V�[��-�T� WҴA�ꜳ��ʑld,��0�n�_ն���E����Aӳ}͂}T�|h��<f�^��Q�uF������l�ů����2�Q�,//�_Wy�?	�w�� ��-#��xTZ��Y��pZK��N��#m�����!�����V����+��00͂<��������l1c�kh���&�Gf3a,6�R�N)��'�0I�Pi�-S.CHW`L-��l�cr�1>�%�no)���o�u+�.r%ev�Ϝ���w��c�������ƶ�4�i�x�@��r���k�f2]�< ��OO��2l��䄳��1�Ƭ�6�
�lA��*�+�M�ܝ�(�19f�"N�{u�Tx��w��16F@Oki�g�3K!L!�d�C�L���P�ViÈ���Q�I�s��3�QN�g�Z��cɨNӴ�)´����x�#��q�Lk���cI��g��Q�uk]92�G ��2�b�h�d$���� (���˳e��Q�
類)�oaTd_Y�D>#&f�"��.�@3���o�00�'f�y����"ژ=��L?V]��)��>�n��h?~��y��y �`�a��& ��)z��r�ro���!m����U�0�_���u�t�����*f��x��0p�6��$��ɹ�SU��Re�CT�a�V���S�5^��uݏ�?~�  ���n��œ��������V����;�׵�ИS�ޣ��1kH�Y�L��L6 �IVZc�d�e�C���B�ź:�H�W�A�Ѯg�h4k�� L�a�0�:��Z[�w�=Ck��ʫ�C��,�3�!�u<�H�ܽ�����1:�Y��F �"����4v��Q��5|�h���k�&Z�/h�p���fQ֘�c�S��H6QK��c]jA�{қƬ�|�� ����G��G�7�c�w��?�q]["J����N���l��1c���������������h���ܸ)����k�*��'���)���:��:C��&�a�h`[c�#PV��$�$sVe�����L��T�&U���0�C�*�bXm3U�� Um�JJ[�52Hzu:��RP�`���?��?~�H�Kc��f���sKe�P��Gdt���>ݔ����f�_9e[�I�S[����h�p��b�:/�	劗uc�n�r�MB��Ώ�4����wųpf�+Ƭ�V��"�?Ķ��
�X�6�����I� ���;y�5Ѳ������c��o�sLG*�0Me�/�P��ǌǌ`fx, naA�rF�*����ɧ�d௖�e�yV�,a
��1�C�M5Ĕx���n�;�iʧ�s��ʅOK��Urq�YhԲ3����0�,�u	Ž�;R�s�8�v�5�ERx�����6�>�c3[�y����-�%�6>n��غ���Ѷя��,�G@M�%	��A��l9� �T3)����� ?�x����3�W
�X$3ߜ�#��������e��u@���:���s�Yd;�1�lc�@�Rz��M�a�P��^cX�QRd��g��F� ��l+�.C��U���}��^��0�xF����|07�XcL�`昙� 3����
˒�KK����4�M���c?��I���&�yofS5��W�b�A<뭤�T���=�w�',eH�߁5�����X,�woQ狸N��~O$�r���l�Yf��k}&7��c�G	C����"7b�ّg(��G(��|VZ�2m ��������n@������W�P����d��grƬS6>##�o�	^�4ժ�&��s͛Nq�ɢ���QPe�I��J�b��56�����2 ��yH{��&f�%�9Tf��A4y�����u�O����ɴ���5�t��>1��c���0�
����ӟ�;�ؗ��f*�X�%�1�Z8*�Eϫ�d���'ccV�by� �P:��_�~������(Bm¥�E�/��:����ф 9��s
�BL�\hi3�2{�B�F�|�w��2���1Z#u���?��
q�9�����!`�����%CpT�(�N*��I��
�긳zj�.��J�Fv&; .�3�N����+E촱{�<���rx�z�lkj�o2�tl�v�6�T�|��p�tj������Ti�UQ�kjSp:�{��@�K}��H;oʞf��|N}7�3j�
�"�$�x#& >���eY��_�'�4�h�&�f-�ɇ�be�	�)��S�6�N�&��
�Z�10�o�N�;��ĠM�ʻ�մ�5m�>��cM�S���/�l	-G�����l�EB.�=v�f5"�����a����1մ{7�(6�g�G�m�HZd�N��q�TnT�v������x��|����mo�|F� ���#�6��������h~%��,ëi����88k��{�=)��)W�CMխ���� �Z�&�����b�r��f�k�'��}��W*��d����1���{L!�,9@����������/e�G�[�\������"{'epk�s�X��1���*n��lܶҘdssN�W
o�j��Ř�=��S_��tDcK�jw�s�3�Z��Yzm��+�X8�O۴�7�8@�m�W��3G���`�60�^�����ƅk��=�L��.�j��e���=���;/YB��#�T��xջ�H�3��].��$��''����ME��z��F{�9�)��>����:���UBm���`Y�:C@DL�%�]X5�!�:L��?�����L�e�J `E��'q4���>;
I�.J9��1��)plJOI�K�͖��ROI��j��h�[��e^�-�����P��4�ޖ:�T�1F|~fǟ[��D��o?~��x�|�2�}�˔r�h�Q��Q9b{��.W ��pH뉌��L�6H����@
�9&�h�4�z-��g���-B'���Y�Mʳ@H������,��o�����}�2�ɵH;T��d��{hف�-������1��O�8�H{��1�v��:�8��hIվ
�>�4!V�[�b��~�,X�eY���5Qdl&5M�{�d�n)=�_��#�@�~��M�̛��<(�#I��
�c�91���Q�^9�M�y^0M)(I?.y=;�[���\�|<)����`a'9�؂:.��'�s��� Rl�h,n�)��F�gm�%FFہ�'���A�G�W$t$�#�.S�!ZY�����xˍ�juU��Vy�>��aG7s� sԪ��%A~˹����u#�)�_��he�Zlm轗�,��&�ԫĨ���C����
�Ԙ��ܧ	����ג���z�v��I[�`c�)����Q��]�k}N��\��:M+P��7����k�S�֖5���	0���g#)k��	�b������U)��)9��6����o?�V `�}q]ۻ3�r;�?�%�ţ���6��B�~YJ}֦�~^m4���> ��H2�����X����;�l���ǌ�>c�3�e��&X�I�10���ӹ�}�����}�/�o�.oI�ܪr���	ɹ�N6��
e��C>*~Y6�N��\uR�*�t2�����Yl���g�����qf���ɣ�L@gS��h��j#a�`�Ψ�~��[aS�bi���:*W?S�E�`�U�������l�Y�a��w&{����j��U�Zv��栖���+��]�2b����֡�|5�I��Z�ۑÍ���-�P�]��<�UH�X{ls� ���'���*l$y�7Zy\Mɨ�@�f<e���[r�lB�]���?�v�a��0?f��x<���/�eI�dӻ%��c��� '�\B��?���{����X�<�ow�&����5]�����i��~��v�]��R����K�-9:�c���cL'�>���QN�����&���/�>�X_�;�c���o��o<s]��Nn�-��~���r��3`�����'�pY�;6��*=P���YY���]�J�� ���l0��]7�#�Ln� P��2[klo�o@��t�\Z��x��Z��� ^��G�]�z�;<�H�
�����@eZm�>S�F�Ik�lB�����!�e����Ә�U���w���3�j��Xg7M�<D� )���g�n�t Xr����Ϭ�+�ʄk�I��4�Ǐ����;��mL�+�^�0����h'7M��Hށ���Ai�{����	�[B	Uٲ���ۏ��oJ�����,���w�Kʈ���a�1��MFm(�,���
i���S�o���I�PcW�>lCKZ��N�>�zF�����m���Y�!��z:�V����?�h@��9��T�=��8��u�&�i[�g�hK%��[���^�:)<���=T�k��i�k�^�#n2�S���}���-1� �\&n�$>.�ǜ�s2�1H������ d�v�����k'�O!C�d��,�`���1�u�$ǟ�A�br���_Af�h���JJ���h^��W����>??q��[pBmBD�{���X���hy}oڿ3ɪ<�a5��F�-���'��|2��FC����O�.��Y �N���q� �i$�������g����W+�F���-��̩�\0  l�{P��w���~��hc�r�Q�j�!�`�ZQ�X���c��d]V��ψ��1���}��m����~bf\�/�We9 A@������"[^��)� <2�����J�?'�K]������C�3H�9����Kf��5{�;� ���ckL9�3�ŵ �1���lt��˦�R��J���>��+�H�/�3&��x����|`�o��|�1�f��>DX��18$[��O�t����m2�J:��Ǥۛ��:���'#e�ܖ�R١���Kʣ��n�>�a�A������׌v]�jEi�pɥ������6�=;����/������ q`��>�!��Jn�S�����$��Tf�]w���C��~�\��yVF�먽@�j�xt�d�Q���B����>�Bd_�4>��S@�E=ό�ޚ�S�k�!�[A|�ߍ�o�t�^d~�Xd��9#ܜ����~�)�.��zw�[򉘦Us|�㑘K��K��~?=~���#�0��Ox��`!�yIK���&m�4��ط	1F|��[�FyO0v�_��n�È�]7�y:���(l�o�L�$Ovѣ��߽?�'l>�匍aylú0��m�i���y��t՗�Xr6D��������;j�i��%�X{"�X�qg��3j����Z�ǯ�T�W
�+��'B2���l<��3
G�0�����m�κ�Y5u5o��,��o#��=&��9Q�s���aR�?�J$� �r_k�R���UBE =�4M��!ǲ� ���?j�W�҇����?3�˲`~<�x,7����-E�1@��kcH�4a�zig���dX˕����g���H�긖�h�,�	t.-��/�E%3&Ę��[i��c���v���L���9����>��ւ�O�g�����}��M���Z��m�S6��������Bzy���1t��� �M/�A>��YUK�Hm��ަ\�iИ2�8��z�cG��k��1��W�V
 ���2lR�Gk��|� I}N�e�i�EZ��� ���Ik[�Z�|�5���$Д�Ej�2b���8��������*�ft�!���� A�~��� ���e^|��Ԝ�H��O I[�G�a��s���tB�2w�1 "�t���|�2�S�2C�Y5"�a'��[	Xj�- �F� ���֤�A�&d*Z���� �C�7j��~�uUέ�$Ɉ7�7M���g�ւ'�K� ��=���V��+?s6Q���Fl���uV,<u���O!M�F&v�S�R��;Z��T��w�?ne1�S�k�W�Cb����1�@{#om�W�>���$��%iy��Ə�����d�a9�x4*=���'1{is ��]��'������oy���P"����	����ei��CH�������ǽ�{"׈=pǁe��B�;�
�g p�c�����XH8@����]-�d,#�^�ʖI���Ӟ���Z�2��^��DX� $��������Ǐ�������?�鏘sb���C������OL�T��ҿ~I�HB�1��c���j��S�����d���	�κ� K�X�m����89�	?D �h� ͎=�d��^i�����H�՘E~h8
V�I�:4�_ڶ�}c�M^ۍ�?�-@��UTs/�3�|� Ƙ�V��w�A3 ���(�=&P�.��Yi�:��S�����w��RZ`��(a�v�&�C���jwj11�V�J�ʧ`�\-��n�A���vP��eC��9���;v`!��B��>����˒�)G���	n�0?f�Z=QR��(�Z�!,9�{fNC�d� �Z�P"���{O�L����1�A3
�"{A��ub�h0e/j�\ISE�k-�y.v#B m�~Ӊg�7-���wuo'�ר��L��'#'P.���|�I1py%�S��Gk�zSÎ��z�+���4ό�V���
����l
�K�%��<̞ ./��}�8l��f�Qz��C�q�Ә|'i��{�k���:��A�'���cHJ� ��[�:���߳�6v���(���;��"|qf��� ��K`2�P1�1�����g�f����i�C)���b���'�����I'~���fm��`/va���[�P�Υ�7��v�Kf�|�HuF�S��yQ��ڏ.�.�<�)�C����g����8y�W�4影�/#"�J�����*���}��YɄ�0�����u���#׹3��������IL��M�/�GD�Z}���Fi������!��PW	�Us%A-���X��R�Ul��0�SJ�!%1��:o��r����~�}y�G�Tߏ�ޯi%�Ja,����</3���BJ��=B��YlA�Pf(i���<ϰ!`��_���� ��@���q�$\�I4�xe�N���B��?p�ݎ=���pJ�W�k�ǳ^qG�KM���m���P�;��.i{(��s�I���j;C9m��������ِ3{�s����Cg�����-�>S��g �^�K���=M[����[�M=��7�gHZkU�Q.�P��[p;�"���`S*K�[rN �2�Rc4Gչ�pP�Y/�z��Q?�*�ZO��v��� ���D��}�Ƭ{W+k�V��]�v��Z�HB�x�� EEۋ�Q��d�o*��ڱ�=Pzh݁���� �Czu�x'����������gzV¼�M�?9�f��1 d63���,�)���M��J������(�����>i�ڕo����1"��X:�XHOjM��3����'��J�:����"�Z��u>1)�;� �]�y��ψ\t΂�i�c^UP;�a�$h���,�f¾R4�̖H�����0�U�� �	k��r͑������ᲕM}t�]7^�&���Tyｿ=��7�����rD4/�u��cc����6l���6N����l�~׉8���~�o1�$��E�Z ��w�S@�%�,��eYV?
�:$�i��~�,{���&S��_��s��#Ĉ�-��y&�:�\��lղ��^;h���j$���Z��m����T,k۫�`O�]��ΊwtW����8\�.z��w���lc+�{�	��;�6�K*�k�Y��J�ju��k�0�+_c)[��Q -ͳ�}��1/7)'ٵ��d[6�����~.[}���!'�Y��=IZ\�},s�! �d�9/nˌ�ܲm�/1;C��0X���ݽ4i�qy��<4����k7S��rr����
r�ڿj��'D���*��6�-ዂ�j���m9���~D�2�\�=Z�Q��O{�=��*�m�ʳ��^Ȣ����V��_e�9�̽�h�klȈ�_{����Ę�,=��j���6��9�ʾ�v�̓aP}���U���'h)�����)�zT����W�0���b�~�C"��a1K�#qW�s�Ζ�v�ۮ�#�1y�S�eJI�k������˘�b4V�췃_��>�IU΂�� ��H6�.� �E���- ��#���ы���"�?�Ґ�hU 01�D�OU!ź2v��>a���H��O�>1d{��Un
Z�0.�
@0-�lt�Vg��cߵ ]�!i��k���8��mO�}�Q�����k��&룹�C�Cb!|��|���[��N�<��W�0DUY��\�ڑ�x����'/i:��w�1��ș%Y'���Ѭ1:1W5pQ{������{�Xӌ�#�O[���=������-��������5�;��5�"+K��/�+`��H���>� �����T�܇�ʸ'�~�~�@����7���z?K�5� M*�v���x�~\J�f�4��m�u��=�1�a��H?!�O�3���~I��˒s��=&0E�3���L��y��>�y�M��K�qG�Iy��]�9�m��*U�1V�£y��2%�� )�e��f���4�G@�$�&�ʺl��d��e��M�(K��;@R��4�O!�����v�ay���A5Cr���|<�#�PPu�'82m����1��>�1%�3ɖIZ#`�RW�6��V��lr�w���*�����{ |DF��������]����wi��!��%@�ϸz-�eŘcR�T��:��cj�����b�U��+f@%ڇv�&��_�D���ھw8�1��y*ac�Y�N��{�eA���2{���@�D'��ɺ?<җ�[@����T{e�Z�}��`j��<fplRk�NP:�6*4a[�8.��4-���Ѥ���՛����z,rp[��\�t�� ��Vu��˘��gU���L�����I�ë{E�Q4��&��r���=G4#�9ˤ���~?rzeϷ���Y��s31��l��^�< A�xQ�>cM������g8y���g�y��,����R��,�����-��Z�P�3EMN�'���L�5��7R����Ȃ��w��8��Sv���E|�Iq�~�"�g�d���>�	�s�x������g�_HZ���#���$�@�V�r抄6�i�0�s:I# i�5R_��P���{B gT�s&����:A� ���<4�
���&��y���ǚ��� f*�)� c��U��=����5�J�p|����3k�W�#��r]���Jj�*�%v`�}� ��2��l��U�`�p&	��� �T��v΍R<i>�<��2DD�/�l\�g
g}��)oz(���jvXr��>�6u��:�V"J-l<��*�V�p�@�$-�|r������ ���j��B�W���/�:�z@S���N��L ؐ]��P;a�s�o,#�#j�#�F娼��Q^��R�_�I���p�tb�����Z��#q$y=TfS�th���f�b�Z�i	�m�y93o�)fɮ��y��Z���-�F���X'[O�� m�}k ���{��3w���N;�>۾�v�Y�ZMC���Y& i�-îӄ_��%`K�� �RF�N�;�ޮ;F"&��U���v������t߲,��ʴƤ��j`mr�Y|��.S��`�Fkl�7	`�����6�8��g�
wƈ~y_�L����5kv��c;g�wn##�N*�x�U-����T�MC�0�2����mzv�֤�/ܫ���g���� �3rt�Hٮ��I��V�A=Sf/��Y{�
LH�zУ\�YڝA%��}�3½�5s	`��'Կژmًji2�� �����4 �/�	�]�d���!��B�_�g@��ؓ))}f��mfs�p�Z��Lg!s<�;H)kʈ�����ڤߩ�`��j,֘�q�7RơD�mf�(���O_C帻� ��g��2��X{��N�G��Yw�wg_�L�J��劼�#B�= ��Lڠ�_Cu����=5�V�v�������z_}�iy"�gg`�@�dma��u��ν�5g�~����x��LJ�����{f�R��R$#��C���_!Ϩv_]?}�:��uL��;�v���H�Ͻu\�zM.ϖa��3������*"l��@J�����'���e.�?/Ӓ�z��Te��?��9�ȷ��B`�0�"]#������WnVZ�I�U�QB:��l<d����W)���s���vB�&~��'�c�샖�����h�벥��J8s�+_���4�P�xy��{C)��2[��Qͫ�QS?��+5d%l<8��Hi�|���Y�`.���UcT��^��wJo}�7G�)��j-���H�
�%�;D{D˱�2�T�1�fS/���}5�0*֚����[���.f�r}?\�[ix�Oᐖ�3}^�ˌ�2�M����_��;���w���M��0&V�6r۫��R2[4����i�r�P^hm�B�Q,y+�ؘ0i��ׅj���E	B��yD4����X��M���������L�S���`�mn��b9e����Xn�ni�Ѻ~�<Md[[��g;�z��MͲP<��PA|<T�#,���� Ӯ�ߎ:��#��Ny�Y�1A�7~|o�ј�e�c�S��e�̽���ky�h�zr5�س���v�~��k��^�Z�YϨ�QhQ]��Y$յ���[!|_��y{��@#�[���9�7v����{ qݏk'"���Eu]K�!z���alL@��w��D���ɹ��0���U��gR�g��˲���O��y���U]�
��1�����������_-r����G÷E���/1�(m� |�M������%oCT�e5maR�h�T���´N����?���W��#��6z{���1w���CT�(S���Jիtz��3��!�N<�}�"�bZk�15��?�m��C������Zp���
��j7A=1�1��&��V�}�>s��쬌�-߅=�Զ3��H`3k3���{��7�=&L�	�������y�����	��!����l��C�k@��e�'	!��8kLu.�c�z2ڦ5%U�hR����ݜ�����}��.��k25��I�:{���k<��^1	4���l�Δc��l�<a�2� z�~i�ǟ����{r����d��^��ݽ:%�ĸ��|�4�c��Jn�.�ߋ��׻١W�Dk1��̹�T���d !3r{��5&����Z�$�� �(V{$�Ȼ�!�X��_L`�YW��$&u���,3�y��1��>1=�n��w�'��J�f�i��d,���=@)<�.2�]Y>kV��T�@`��'Ɉ�����z��yDB��c,��a�f�^�̖���C��Z��:���l�
�M�*/3m�	H���.���)�rHΖUKX۶q<RO�i�c$dNb�,"/���y�i�&�K��C��x�l�(��e8{iIH�g�C��x������ �|�t���1�̥��$��4�&.�d�Z&0\^�>^�\[��w��x�����3�#�:̵�uO��ny�q���)�)u$g1˞<�`LV���E�#,Ym�m2�e��g,a�ݻ���&�����:��P��h�(9҉�M�d)���#����Y�ZX��w�'�4����mW�����vr�R}��8@�L��c��Ǉ��T�י��Ө�hh3�-&�X��׸l-ዯ����gm&[� ��ϰ��Zu�֬�\a0�1������T���i*��_){�=�Z�18,B�1�0���l@��YcJ�%���>�ek+/yՙ����!+�<�2�>��2Q����*P5"r���7�|�z`e��sE{�:��c�m{����i\���Y��71f\s±ʳS^p�@���i[�1V���7k��G"��}g�i�1��y���?�9�,2�l� &Xxq3T�(�Q�&��cv
�&�e�Y��s�����ۄ���L�Yg��@g�\�E��UR��33Ƙ����J�9[X��b?J���چpp2\#30fp�dc�9wuPCXH �r*�Ӕ��/f�/���[����-d����Z�ܽz�j��l��= ������˶i��7�g�+x�hV;L>&�����E��F��L*�c���K�eĆD�M�	���g	ꁅ�գ����t{���r�=,}�{����� )=P~��������MS�5.I�^�j�}F��*y1?�s���K*I�hR��e>x8���a>�~Z̷O|�&�n�pΥ�m�,T����2��d�#E�O)��S�Oӭ���2z�b����ܸh������_����@mWyR��2 ���\k���ԦޢԺ��DZ{��3��w>z�?*{���+�M62�� �{`�����G�l.��s����w����<(>�3�<����h�{�e���	0�����d�IJ���k�ٸ�\c$?�J�Ⱜ�~kmEf}�$l��R�=)�$hg��kB�Q?G��� "ǨH�n�A&������2�(sӔ�ev�5����I^��"(�@���|�^Z<�cX���q-�%����B�ݬ�A�_.9��ə�����83���9#��O��ŷ��Շ!l�� lbnj���򡶍6z��*�~Ɇ�=߈��Y�`J�w>}vd�i1Wrc-Y8zq��&&��+6]
��m�d��]7|�m8V�:Z�5�!��LL&>{�{$wzQ�g�6�{�g,�}�����P�ه�9���>ߨ>�,8��ֹ�C�Q!f�ڴ?#ڳI�����H��}�{�v?��S��Y�����k�W���A��"�9Gk�	06��a`B��,˜U�!��)%` �~yy��ȷQ�����2Ɓ,&B��f��[�f�bf2�|||`������ۏ�
�4lp/��%��vګ�XYH�q~7�&i9�$�bzu��@��8��Z��)�Ulr��Ɵ[��*��y8j@�_����B�V־��Ռ�,����T6w��k[e�A�rN-ֳ����
��Y%M����<�ǩ���[��/���2u�{�j
o�M��4�1[ܶT%D9�#{�>-̏|F`�2'�J�ǅ���[��͕�>*{�Hԁ�C����Ly�k�C�g�=(���6j���vρ쨹����%ؚ�Z��S��� Vƍ?��˓14{`�/�'�spqdu9�0/3�)P�~��1��1Ͽ�x<
^�8�1z���6}���%. �lYV�,�Dx}LB��E��!g�1�v�c�Y���,� �f��J����+�	�#�Nr��^P������Gtm&�]C�@//-�5c�˾��ɼ�s�V1��8�q�� �����Fy��4�]�#�b�fec4}U��c�0._�v���eQ��2X� m\v0�&�{�P<����砅FB5�5<WO��`:�e��[.9��#���3rN�Ů�����'M	��M<юM6�Y{�k�v��%ˡ��:$�=�~�ZCu�u�o�uVZc�@L��㶠S#L8�l�T"9�ܤ��^vT�wٿ��ؾiL��vK������09�cIvbL䘉�9�M�7!9	���+�X
���1XX3�O�m�<͘n��?5���&������p �a�9"���˥�/bth�?V�]�Hi}>*�z@[/u��s#��N�GD[������[�a�=�{M�2Ҧ�g�'���T'g05u�QU����H��M|F�<Y	c�׆�)�B貈�]��Cϫ�ǆQƕ�Hʯ�y�`q\j�F/�[F=�����[Z׿8�~O{qU{8����Ɋ���#�$������0�er"<�up��Y�l*+�K�#�}E=���G�f"�`�m bvz��2�M��}�H�cb8��	�� k���^yNޮ.?2�l�͈GDz\i�Q����mUX����j�M)�~R�`����#�����㣺~������H�}�v�i�R4P�U�YZj���̉�Q�>_d��LSJ'԰��(^�-o���|�@��s���
�*M(�N�SFr��~8=�n�9�*���H���[�U��b�5F�ݖ�c�~Z�h��J=�Y?�d�ʼ�_��񿥭{��i1�n���[�.ƈ��^Tȼ^٦�ѯ��l�)m�+���:��P?���'��_�,9�� F$���Đ������&��S4�Lv����� :[�M�,��Æ�F&з�[@�<�X���P��ѬW5K8�bW�.��F�G����*;w��յ�����W�(�q�"3G ̭�v�\�7�>=wHGֲH�Ŗ ~/��ܻg�?f��|�Yԥ)����	\-��4��=�d�Lי|H�b�r� �H��a�C����˲��Tʕ^�g�֯3��w&ãN�7��bl�?+G��wGjAb^#�{�H��3���n�O�h��W�K��Pn]O�����&���W�sH3b�w��?��4�Mw6>�5J{��d@Q�w��Bu=�c��sr0�ǌ�/s(1�I���ᗔ��g?�,	0�XT��L0��~�~&�H69�$�1DD$0L���O&~>�\�=�)��Ȕ��-�1���!{G%���7�� ���!�0h�'�2�n;��8OS�%��ԃ-�x<B36% ��B�U�A�����*RKZ��U,�;��@��F���/�9P�n�����V��{!od��#�I�]�����8��{�A����ѾW1��D�Ne��k�����rO�9��w�jg�T���z��s�6vS'#}�a�����Ƈm������F֍#c����r$�������{~����M�z���٤�2�%՝A�P���i��J��8�΅��i�OQoL�����X���&��D�!���   ؔ�;,)JN�_�kD�2o�;�i������垖��1�jU��l~'��1)l���������,Ӛ�F��d�����Fw�&��ʹZ��3eQ���S�R��:�kG�UB�y�R��J��'�M~�DS��Ȇ�m��<R^���|�24������	׀���7�z��y	[��R^��ƣ6�g�m�	�1�Mb�K�+�i��Lp
�cY����Z�3F=]3���8`�4&�~���,KX�K����_��l%3�
1��A	UD���f�!�4�/ �f�c crXF��-���Z��/��>?g�i~���	y�4�E,�]������D��kd�:lh:��j�`WS�w3o�=�ʊ�l�>�@�2r��hDmJ�F1�z[l ��_�t���ZD_	4ϔ�c+F�%ؔ�9�yF���
�ɳ6U����P����@���1�{"C'�����)���� 6��du�.�ߵ~�YKi�dE��h���nHd?	|~��!Y�C��=�7��b#z�|վ�
$Iă��H3.�Ln^%䞱�R{�fZ�=͙5�ߞ��6˔���Z��(����7Y��H� �	�f~_Ddfe��O��8'9�\7��p��g$��y��լ��x���� �@T ����yt>�����T�PU�|��_a)�o}��l�h*�ӟň� P�i�@��'Z�C�uE��]��r�C�,/��z������?�K-*)��̬!���@IT|��.���h�t?�-r|3��)n�#3E[IC�H�3��`v���~�сF'#��\QM����u@�m��V�-�T����7�3�}�� �$(��Yl/J�'6�^�>k1��=10�S�@d0�9�:�!�:�t;�g��]�E[���GQ��=��n �`*G��k5
L��NZ��X���'Rs����y�Oc��#o]�S�.��kK��gՈ�sU^�?��&hg��˶����ܛ{��{���q/��U�-��2�[�����7�>����X]u�i�j_K)�!{vҊAHqo:�XJ��Qp��r�wkH)b��\���qUJ�K�����[�'�J͍����R�:GE)*��+&�\1�D�	�ʟ�\1�@X�ú������/KS\�;�kR 	l/�%��}H)e晉G��-���C}$T?ۆ��R�s �rh|,5h�b��6�p���o�g6�fR������Al�G������� ���(�#9[���%Α}�1�};��C��ֹo܇Q	L����l�Qڽ���G���g��z�\�l�t���W��S�$L'�ۻz�?�lp��^���Y��T���D�ӌ�Ѧ7������ETsff3;@�fB���2�B�p>���;��q���*yY�r`�,5ɺ��="3�g?�-Pڿ4Y&���I6�58��|�I�����3�l���4��%%�}P�R^����g��q�Y&��v-6�+�Q�iI����̳� �� a~=`��$���֡fх��}f��3�*�)��|f�h�W���M��:zggA�Y&O�5��WͯV��4u��"2�C�<_y���<3�ez?++��j��o����U�����.�B	����)�g����@.�!!�P�Ae��w1�b
���"qV��"D��WXi��v��r{ؽ���R�i�H��y2��# ��BY�\:g�YJ8�|�k�m���Vz�{4��i�(S�!D\.K�2�w������64c�</Ŝ<c#�R.��/���޹6M��^�YHi@��Jޓ��p8�d�{��>�<�_̴��M`�ˁ�\S6�v�������%���0�=��|be�蝦���Ky�j���ؙ�;y2�!6���d��=C,2B���d���Y��ߍ����Jfe��r��C�@i�d�sR5�۩����f���2�ތ�W�st�~yJ).��n��bY�s����[)��7�����c"�
&SJ�(&(契�6
@,�*WVs-�ٿiY��3�,x�f�1��A�+���̰��I�&6���mZِºH�[�WJɬK��{0�;�{�W�ޏ����է���wa�s���Ov`v��麧��n��"t��{��P@A��r?u5�����U���'ҏ�Q��,�u���(E�S�䜕SJ�����W& ��JĜ�W��\�)#_H����գ����N��,�qOzk�H��bY Fs�".,����v�'���>:�!�����7�B��������r�r��||(��b����Y�+J)�S!Rb���bDt�PNp��W�1'k�޽wo���L�� 	�g3v�DqFEK��	�/�9a�n�w}��͔`��&�ߋI��������vIH�Xp���]j���G�&��zԋū���������Q�������~�VD�J��X��+��@���f(˜?ø��Ѧ[�s�EҪ���,t���r�H�Ɨmb<%C����@�uGG���X��1��;����= �E-=������ɖD�!y���;��"R(���BD9�9W��)�\���Xff4��dL ��%Ęקln��Ō�� ��Y;� r�I��_����0�D��yP�Mdi�&���*������}6#����enL��b>c����}3-p����Ig�3A��&���<�B���N2�D� M�<�͏�:͙��\��}��2�Q�^z�ϐ�5z�ͽ�|d ��_�3\C�p7��6�-c9W}o��Ȳrf��j_ș~<����,�i���y�"�������b(�e��=�h]��H�m��Öm%#ʷ��#��-�g�D� ��
LbV�B���-� ��@�쟉H�)� ��&����KA�f2ፀ��,�6��r�(�-T�`D�����1���{&�ƌ�`�y���07p.K��S9V��L)�j��s���<ٮe��-�=�O�� ���d_�ʣ`��f7
+b�r[�m0���Ȅ{�(]1* X�����gI���8KJ)W��>�m�ݗs$c�
Lv%�2�0��ڟ0��s~OM$3?������:򈜵���{D�ӯ�=Y}�>���gM)�m^��hۛt��q�L���c��R��eo�%�Ĺ4%^�T����J�`�&iOG2�M	`�!1Y&-����t��1D�%U��w�����"n�~��C��.����� ������-/���[�L��n���ou5�?�z�˥lDT�d���6�Y�M4�V�2]@6��a�mZ��$���N���%��y.gR1�Z�����G��N�bz��cg�>}�Q?�fu����L[yqk��R��l裈m3p�s����MI��s��g+����|w9.yC�����R��ׯ:��M�S`k��p������U R�WM~/#��{�}sEΥ�=��b)ERy9�=��w.ߓ��|���#P�bl���g���m�#?w�m�A���u���)�3}����;�{����X�G�Q�l���J�FJ�S���< �1ᖲc�$�r�Jwq�r$9��e�"^ֿE� ��r-s�� �x�kVt�{�5^���
PM��- ����)3�1������d쎘. S�9q�\p��7��6;W��D,���Dd��9O�(����{��'�∺U�6��e޲����w�W��h�� 4��"�;w���2�Z�b�7뫤aN�A���<.�&���G��?Ȓ�מ*�xY������<�\�ʍe-�.zm�ϓ���N�\�����Ϛx�2��<��[O���2[B2"u���=��VPн��+A�3d��k@O�ޏX�G,'z�ׄ���u��Ԛ�G}aVr5��I�^�矱Ng���w2Խ?ϟ�^(��%n��5�2�.W�+ACr�H�88\
A�8�B�J�P-Pr�.73��,���2P,�LP$P,�%Êo�1��O�H�9#՜VfȪ�n|���d���u������o=ï�]�7��Ȍ`��#�ǚ&��#&��Џ3���Y�\~1F�/�2c2�Gx�u#�O2�͹�SG!���Q	�
�:�Z*I:���'iw���_9�3:�4¤��,Ki�gS,�n��e�H}->�
�>��	�����wuF�{��RN �	���Q��yg�h��st�x��G\t����!�L�
r~S)5{ٙ1�3�L�'|:g$�w��X��\����&� �Bt9r @�jW�έb ��L�Ѻ".bX�ۏ�r��?Q��|�0���f�k�:����J��ϔ���qiJ]Ih�7�ՂvmN,f)���M��<O��"�ͮ#O�M�a���4��gi�<����5)�ڹV��=��ԛ8�1���cA-���޵>Ѽ� �;�k�	���˥-�\���/�ݼ�	f��l� }����	�k���<�����[�лs�䧩��ϻ9�@����D*�3
����^?d�3�w���L�S�/	�9�1�*cڕ`+%�#	��x��b�n[�)�r��5 VE���7�J��) ������r8e��*  �P���s��P܎�o&BI�\:z�e����	�w2��i�r2�l�_�K��\����=.˂��Ҙյ	����dͩ�ٜ����q�2��������π�'���H`���vG�?탒��X2jO�/k�uA��r�}ʦ��~��rdFmR줽� �����iW��r�5��o�e���>`H�p�������㈢JӀɵd�������h�zf�%V���=XF"�w�9a�=:��3�@�i����^��92�u���Z��<�7�/�ge�/��X����̹�/����eOȏ?��j�k�RU�5ϥu��r[��sooo "���1 ��8���G�O�˂e�5����<����\v� O��i�P�D9]QL	�Ϧ�s*�"B�!�6o�w��[�y$[B��ɏ�'�_<���du��p}]�p.���?�I�&6��d5�&G��v��a9,a��Lg�գ��3�#yh�%ڙl-s �k"��:v��{+�X=���>Ja�9[��;�[��k�^�q���������`ɈQ=�?hI��"X�0���oV���I3�>\?*��$-=�6�nt$�����;˺�Hm��>�wR̊�����]�o��g+A�	뺶V�c|O\�[2��C.���xN��g�H%�<& �R�<?�e]E	h���x�W%c�`,פ�1&W��:?�P���қ�/9���vY	�Y��o'�#�Lsw�� �H�������ڸ��O��I�h^i/,a�򌒉���=;׉�������!���t]������^��^�����6G���%+�F��Y��_����BW���2�R,&��~�:hλSY<���� �g��Z��
,j��������
u5� �ܑq@��zݖui���9�e�e���(��.� 8�U%,.m��23��5�ru�I%��Zp'aM+��g �3�\.W\�o_���k����
	k@+>>>@Dx���n�B�^�X����3�b3����41IT����Â<K4�|xΘ��vi��=*g6��T��
�9�(��I`R�D*"�+h��,2�����f|y�^~<ݧ
�Ez"N�4
�����1��Ca
g��l[�s�|c4����)M�˭d�ѹ��8{>K7O����T�u���`�x���2'���w��ne�C*/C�#c���w�z���ofU
;}���{7�o�uw{$O�H���B����BX�˲�z���ǂ��Y�/f��� &�+��x��
�L)�  !��Hٖ^-)n~�.W\.����)�I���b�G����;1F��0ǥ<�=!�L>�R�'�RD��#�B\A.�/���7\�Wx�4�N�OYr��D�3�Y���4�ю�^��ɥ�um`n�]X������L�~S�vz}��Y����g޹e��R��	&6���O^O�֔����o�N�[:���X��y;VS�Ms<�6�d�ԥ�)x�9�k�w��AV=�Q�<�Kޗ�m�iҲ�y+{@PJ/;�NĮ���yF�#����ǩ�l~w���W�}|��<����{�s�9RBy���V�^�o���=�@�|���݊?�`P���Y_e����L%�1EJ �#!���?�D��	��_������W��������+n�� 5@ʿ���+6��sw���h�T?Lձ�?��P�Q����χ��>�,?KbL�5�gϓ�9L�YI)f����˛BL�i,pH~(�>rO����i��M���ɍBF8[����D�6`�M��XLF��6�u]��0`={	�h0��{ɢ��� !)���0��R4��q6��i�Ǵ}�Ӿ�I�2�5��sL�� ����5O*�2��=���������Kn�2�1V�����e��Z�u>[ҀLv�4DT����j�Φc�"�B��o�>'��:�-�c7��+b��^��^��Xޱz��e��mi��Y�D�0I��g"R	���3!g�)����_�{�2�鼃,ۨEja֠N)���N+ym�\ϗ)^���.��g�N�C��4�N:N�~dv�����2 7����W�K��y�1
g��|�2bM{��Le^��nò�/��,����(E�*'���6l�����7�gE��̫��Z�
��g�#<"���8�%�����s�JJD���A�WOv�E���}�)�P�g�c������k�*u�q$�a���4��ئoYpd[��2���(ͻ���������Y�݅�SE�l9]ṙ��4Y�֫�P��$�d� *���蘒����_��,y��<qf�-Z�En�Ψ ����S��f���В�9m�+s��2�f �l_����Y���\���% ?;�7������<���\��
|Y�������qd2�i_��ٞ#�9���Q݈������r���=��[��|$V"v)V��}��z�Hf������
��~��4aY�Z���UpM����T�-K���3�0���r^I�})�\ ��|�~�{���iS�x�2��]\2)���;HN${R���H�B�c BXkv�6��V��ZMץFd�9�b�D����.��֨ ����!E EdD�b���-/�k���Y��'+�L�[���G������ɠ}�F`�����w�{,{Qo�mޕ}p����x1a�������f2z����lsL���q�k��R@P2����)�+ �eA(�ᑉE慴|3a끎���������{��
T���Κ���+󵦔�Hx�-��5��$���	�xKj�$���z��f^��cԄ����YfvK���0�����HEY��'���}p��]��,M�3پ�m��V?���{��3�~Z������h�����rOHN)!��1� �s�1`+ޖ�r���.���,��t]<~�|�2K�@�@�T�bBMc$ >կ2�%�g���u��vy6�'G���"~`��{�p��8Q3��R7�ɴ�o��`z�]��0������������x�Rz�(���fw��)��
����>� �^��wP�`Vk��6�z&����h�y?�����'��i0]3>�g�H��@Ϩ?_�Y�m$����c��������X�3U�k���m���g�n.(�-������g�J�u���e�'(�?_)9P��yD���c--�M�Ņ %Ą�S\�DMH�\�@1*���u���̉��)�m\c�~����Ǟ�s�% S���D&d�A|��3)rR8G�6��#�ُ��_Ê5�goaZ���ҧI��<��*F� zkL%��Ծ�Z�x<�y������(���X��֌� ��T,�H��U�X���&��Ϫ �h^�{��9
h����k �>��J$ŘԌ��&�/[�g*ƍ"6r)�s�U�qAI� ���gԿ޹�-�%X����F�~��� �E���Q
���: ����Џ�[, 5 ���Ϝx=E�{��R}9�\d8���N��I��dF=��AnEּ�~+:�5Lfa!%%$��(�2���Y�ih�ާTޖ:��1����4�i��ה��j������!1�c+����c��Ӡg���&G�jZ��ŕM�f��#��OͲxV��0���{�{�\��O��מ�����VS6g6�0�7Q�1���TB��h~�����_��;���M��l�M`�~���^��`h�ó���#�ٙkk���B�-��m�[�Ȗ�����|2��o�3���0���\��}��3r'`�1�|_J!�i��o������;+�f�x��'�9&����"/�������#�����D	4��V{�),W��_��X����e�9&x"����*mf@_���r��z��rm"l]e@y0�n7�fz��<`�h�7�����XLل���I��וb�I~���a�y��㜫P���E�X�,�H�1��d��kM���@3!�i��9 ����l,L�$]>��}�~�
.˲l�����qc'��Tޗw�r���{kR-�*�������c�����=�P���W����;�8��;����wLD�����{�gϬ.�V{���ϥ�^ې�*��#����gw7���"���9�k�TZJ�>��a��=(��#�����ֲ#0�YN�,{׵�KO����޺G��XF��^/Ş�u:@.Si��\��a��r�2�)%���2~s��Jj���_� �"���bʬ&w�a��$JTP�7�l��BN���906q�J���5)���@6����ɠ�	SJ��i�)$�sF�Rڢ�8 H�D�y�||z��4������h�ӥ.���Ӭ��w~o������t;�q��H���L�`�����)S���^e�:f���q���ɠR�728�6s�:�a�k��m��t����RR��#,`J��0�?ߘR�V鹿7��^+�R��{�������.Gm|պp��v@�h��/��C����>�g>G}�nX\��8�#��L���k�����-�V��-��ڍ�W@�\·��s3�,�$ρ@��l�WB�Sv�}+D��O�N�LyY��UD#69���M�O���''�s�3���R��K4^�N�0c@v��ri�ԽXO�!�e3`���gFV��H��5i`?j�+7f�i���zVx6�c�8��u��ƌ����2�{į2�T}Ru�����پ^G�tO��	�!K(�#�����|��T�9�^����;]<�F|��<�=�����P��
�.o�L[���h��1��6�cg�^�W���u�y<��7&�)������-%�ۀ.��͘2{S�4�P�/�q�U}�m�3Ʌ-'�s.���~�	���2��_d1c	�¥��굵�+�a'�<��:�:��L�=Sg-8ۄf�P�7��=A�J��P�!�]�9b�83M� M/N#s�W�+R�hV�>��d������$�Oz�55��K׳�3�I�}��Ks;����<i��]K�w��7����;�(�TTk�%=3�g����f�Ӿl�=}�s��=!��,Sʋ� W�r�7�/��3���gZ���������V�{ٞ�,�LJ 9���=a�1�CJ7�YH};�T/�%���R>�6�Bb���컉Psl�wooo�;����yY.UsZ�B,>K�g09w��I5a�1��o�\.H)���d�/l�#x�`Y<�_�Rl6y��o�|�h�����h�-�뷱��T;��,�&�<};t�9���l2���m�ٰ�`i�"�gn}�9��g(�||�bQ�!ڧh�����0�RcD̙g#���N0�H��ll�s4�y(�]�,굃���[��h�0c+�]*'��=���0D�Y�׮���;fE�B�����7/�{�����/��)a)�Y�d������������[�\u"3�V���DZ̀Z1��5�x��6?�X��Pr[�sGV��98�.�~��xĘ뗯! ����Ɇ5`Sk ��zmm�
"f4#R9cA��`ʏ�% sY��x�õ�y �?_�>����JUF��s~W6��>w�;�pl��f�Ti��'
='ך�d�uRs��u�� �3̿g����X��D+C��3�bI������g+��J$�Ӌ���E��ՕeKe?f�����X9�e��J	s$g�	����[O�R�@�h�0�	 f�Eu�sy}�3���/��{�1C�ۥ�Kጩ�R��5cM�I+��TLB�g�/���#��JJ6���\�)�]�Ŕ���K�T �Ka� e�-% A�C�_&�B��ǋ��;�K@���ȃ��٠-'��|�c���}/�6w�uk�Z�[�8J��N���>1�;����F؁@�ޑ)%�/"��19�VNE�z$@�=�3��%���$jX��V�9jߙy63%�ذ�q�.h�����2u�8��Y��c�O:�ܿ�c�D��EO}�m��L��w�D���*�u��嘨خ^�ɜ�2�r�饶�Q����:��� +�08�U0�dFIw�fH���/���������Q>���x�|%�Zʲ~�R�@����y�T��a�)�d�. ��X�i� F�ₗ �QB1���?�/�D��7��p��z���&O&�e��R�Р��Upޒl���萺���v��J4���I� ځF1q�E.�s���ϋ3��g	��u�X���ń9�syd��.r#�,�xFF��2���
!Tד�:���M[�$�-�mY��AN�N��Nt,��� G�Kv>��Ba��Ԋ��Ig���;�����
���,�?���Osok�6a/_U�]h�_�-��]����=���r����9G��)�˗Y���v�"q�9Iis��	�0��jɜ#/V-�<�R�<�PI��
�)O(��y?N�}��d��� )D����7��X�9Aj5'�<,]�=�����\&��1% gAu��Y�rt9 x�4@�oI�]4�zL�j�Z��$����m�֟J���&TIL�'�ۭ��)�s�-�Tb���a�F�R^S��w�%�.ν��˴�|�������i�c�;V����F�X�����tY#�"�u�	�_^b6� �jVE����yN�̓l�ղ�|�� �y�e �h���Q���|	S������4J���m<�C;��w.�emy�ϼރ��"ԏր�k��g ��f$,]Gyc-�:�����ʵ����x�����}h cڛ�G�F�b9���Xo���-����Rz���NuO��h3�m0j���@�&$*9-R
��T2τ��E1>���r�aE��\b�ϘqNX���9 )Du�'	(��˧)�rlɦ�������g�k�����������7|�re����Ҁ�	�:��fӰX�r����x�e�Jj��5e�����O`"�Y��ϊ	��Y�j> xq���rB���w����I�I	9��4�Lz����tj�:�gah2,�{�>ì{�������2�n��@��������^�ǵ'�`��`u�,�'�_��L�L�����S"i�g}'ed�"�1�=��=j��� L���N���{%83����\���_yY.��P�kfvK��X@&ag2tY�bS�#n��^�E ��ۿ�?���}��_`�ci�ٹ7�����FOm�̶��q��543��n-�;v('�2�o�]�/�<��c&�,d4Tf�{Ē���U�<�#s�3��g�R�E�K(��oe�Wkm?Q�]Od���[T�'>꽇^�AW
����)���&mb|������-��4�ϔ#F�w|þu�~��^��/�����wx�D�dtXS�i΃S�4[?ӎ���lq5�u��7f۔F����Ӳ�L��:C?�PL�{���;�ϖ�<��'������8�by	��_���7���7������@�2]��H��Jj�)aY.9��gp)S���3�T�������:/�Q����v���R0Hsb�g����s���8�A<kN��La�����X��2�?z���&7�{S�h��^�٧�h��d�NBn�u���ɦJ p��t�2�e&Bޒ3�F5{���U�w����M^���1�:J^b���g+��?,�}M=΁c��g��J'��;�V	�}�р��[�q �>ڄ p��5SvP�m% 	pA�	H�Iڷ�R�e�opDxw?�}k�K@�����������������h-V�L���(�ǽ�	�CD�	J�s=�9���?by��:��{���U�HJi�}Ĕ�r�Z$-/k��Lk3'��pŴ����,����$��������>��S�M���l_����fAYO,8fx���DnP����L����=&G3La�,[l[��=zA4ֵ�5{�b�2�MF��Yy9�O>^�Cd��y*�$��f����c&e���|_����k̈��̯���`j��L�Z�e0{�P�%rL8�%�^Z9z�h�;�ס�
ZEj�� ��~o�����Y��9����~_�Hu�����@n.�ާ\b�eYviƤ��q�Hͭ�t,�c�I��b���b[��l.��sW�2SJ�����-��/�������?����.H��\�۞��r�M�︬�⽈�>���`�1#T)��$8#��H�<�7� ��kf��R�Z�%��Wi��d�Nf]�J3!��+���n_���q�S'����T�Ǩ��2��(�#��/����4C��h��%`F��" �	���̩�����>S��������] �g��/�C
X�XDE9R�X���wM�����J����u-�V٫S,X�P�c�u�b�J���kp#�2��~�/������7�5!|l��#��d&�y˖˥nw-~�vs�d�s\Z∆�t֬ݰ�΁�|�G�ce�m`�Y�s?S��؞�V��.�V��Ľ6�l{�!����{�N9Q��V3�.�U���fn)�wy��9+ҝD~�v�e5�ꎵ�̽�5����w.�,�X{>S��_*�]2<c~�<��H�yIK�Cy~�:����JqDH��r#�r��	ӳ�e  �>��#�S,�Z������K�ؔ>}�s������� r�����`���9M>S�lJG�KT�f�{!,��m�Z��7�p��{��g����(P!iJ��]'@��t�=�C�H��{�LF�92]r�����MMW��	�u�|����3�k�J��g��T�x������ID#s��H�椽ٺ\{./3��=�G����5��9�jT��Ӧq��o�9�X��\<���z���Q������T�
F���I�5��l|�+���I�V ��L���q���(�`ʲ��L���bs;�d�\. �u}B��$�J]�,뺂��c�@�����"�� �5'	S,y�6���'J�����`�^+ �K�M��OK��ʿ�?)КQ�jνC�d�|�:�O����d�(97f��P1�s7�>Z��tf1�ܭ���\�\��h�!�����4��<C��!?���<�/=9�ֵ��2�b�t�9ז�����܇�<�sTЁ5�/r�Ԍ�~�\��(9��^�K٧3ʀ|�ݬX����ȝ����(�׾��Ak-�~��7z0G�To��<����3��9b�A�Gb��Y
g�����������F�r�U`<������G$��E�\�+�x��z�`Y,���z����zLV��s�4�pH1�٤T�e8�'�>3-ɦ����R���,��#�7��/�@~��<S �����n����Dmp�J�x���eY
�M��j�������`������ԔH���MU����5xɊZ ���E�9V���s�����7VT�sͰ��с*3m?*��DfYL�X	?�QR���Z�t �!�� ���v���q������:�i�����}��S���YP����S������$���h��Y���j��q`5���iB�
O�L�T��g 8���F�ނ���܄3�&�X�MV�Up:BG9 �;_]�����G>�$;��d��0~�λ�%?��s2�B��q*`*� 
T4����g�����~��XO��Nߠ5W	zdP�dm���g��gi�����I���|��}�3PT��~ւ�թg�쀻b���Q�:jF��ƭ\��t��ZI�G��f���j+��`�;K?�{Yn>SzJPT,���2��Zp���ϱ�Gi�4|��<�&�#�A�j�c(8!����'���i�J��ܛ�{�QF9��f@'a&��'�;Gy�^��s7��?�Y�'�v����B_�j�!��io.�i_^�Q�,It�J�YXEn�'U�<��I�t�/�"�����Z��{�	��`?���C����Q��e^���gJ�a�u?���b2X�Y��(���z���A���TD�R4�+���{cњG<f�������~����y���|����ۃ>���3>gdWqhr��f�W(�rm�cI����p)!�֭��~�:ҥ�к���l��c	���?���g���9�r� ��� ��CHp����:"�GY�M"�x����X��&����i<��N䊹�ˮ��O�H���O�q��&�R�����|���Q��Q#��m�����)�%��2��L�Q��y��l�;ˬᜫ%6��eu���&}�Ѣ+�g}�3@�壤��Y���Q���/b�����nTҜo���0�{ӥ��9R������9��V�+ T	���e�x�n�M�$�E�7~u=s��lm��ϣ������T�>������h��G�3��[眽G��l�s��x���J]f��L9R�G��qy����K"B�ME�
H�Eo�6!��bF��}0�����ǰ}/����V�e�D���%�
��g��H r 9�B�����
���y�}�lR�T�E��d6�h�#u�^R:&��� -�����V��r� 1���I#}w�pT}!�z!��rSG�bj�47�n��X��Wcr�	���kW�u.�b,9���ؙ՝�.�|̬/�t%!y��'��|&��%���nb��c	�j�%�Q�Ŭ����dߝ����(�A2��o}}�L���}�3��]���ײv`V' �IP��k1U~�frOА~6̼sߣ7��)ɽײ棔Y�W���Ǖ�GD�C�[�q���uY���y\�Mi�_W��s�A�lrk��>�OeO�k�z�ۃ��0��$��/���H�����u��a]3ؽ,K��-źU��J6/����H9�}"`u8#r�O�y��(� �1���0r�<��A��T뱴/n�Z �������%�L�yɨ�*OH��i�^�f�G7�g0p/2�O,rZ�
�m63 )��jE_1�U �3L�����>c1K�g=�!��G�ӝ�}�^��g�T~R��=�[י��+��)s�����=����E,����QS5��V���YfƉ�`����4�.+��_�:U��t�Xu/��23�`��@0���C~V�߲5���2��W��t�~玲�_+/� !��Z �NtF�I�'K--�<#	�7`�F�_�K��w+�Y�5�^~A�JP��~j����9)�rje����m*�r�l�9�--���#��L��$�=��Gk|r��Ͼ��g��Y�,)G�˖��s�;k�jy�ٲo$ |�SB�����{~eK��̸�{���櫙BK48{e��\���;|f���g����[�="��^.׸� I)!��E/�m�װ�K�N���+R�)֍�f.�]8�̟Z4\iТx�fo�.�s�˨�%`a��V�<Y�/<��߂�Hpl�sD��!��{Ĵf�[�ܙqEr���J��!+�zH���ŔaK 0�m�GbaU�~"_}�(Qa~�{5��d��� u��e�|�@匘Zi�e��4�E��\�����3�!AGOtE�z��T�c�<<X��Li%$���;��n�x+S��6��#9t�F&�^N���-%��i��s�Ɨ�'�/`��g&�D,�h��JB�e.���6����X�'�c*��Gʈ|g����Yx��^9����Z��| ra4���[_�ߚ���O�6��v��y���r�7�es�b�A8	p�!��pɁ"@�@H��Kr����ѵ 3�� �!���K��X��6LI�m-83���$�}��שg�K@f`�7��P�3�Y�9�*�G�F��cy�(�"�s���-�p6rn�/�Y,z��t��5�֌�.��)�zڬ�������N�%:j�H)0�'EȞ�.%+7c-���*3�D�S+����;��7�?(>"ֺ��`��_!�n���|Gw!M6�\Ȭ�Gm��z`S�i�R�Ĳ�9��5?�UDʰ�q�z��XSm豆	��D2# OXhA�V�#ŀ	q]�.�u���S^c.q+�ð���@�a3z��	izX�s5S��ϩ�j�����)�&-�d.�:'��Y��pD��L)=�xh�)P�R,F�?׾o���J���b���3��P�s�ܨ�	��#�L��凫�֌���ޓ�`zɽ�f��N)>P�znH���2��I����`��n�75K� h�$��0�Z��&�k� 'e	K��8���.�6(��&d����ws���zy8���8�{���n���9��娜f*�R�;��K��-K�NÑ�F�}��?�`���0��r��v�ޟڈ-�S��)??=y^�(�����}���̤�Wf"t�T�;Lȥ�߭���X�.����TU�~�k���T2�?o�_�t��ƣ��g�ߋ��<�8b$��=�wOF�|���D�Sh�`�H�/s3U?Q("�o(�b���Hp �Ņ������V�倫JR����}��.�� ˲T�X��j{���r�8EK���<�������ˏ�z��5��<��g���0�����G�������>�è�~���Q`̢���~D�m}��{$۱X��"'�f�yTA���<#���A�\�@��Q�f�Հ>[�����1��۔~�� ���Q��Q9�#د�9�\�������g��Pny��hb��U��{}�����Ϣ�efţ绩+}�KH��Y��z�@q��G��3cE���z��Գ2��+����w��qgXl�g�~;�j.��s%����f��Έ�'D9G7Q����+�@p)餘r�j�,�$e���/G�y��S�����g�s�����B�3��p�'3�Pr�c��gV- y�����f���#��p.��h�^������X-��rwڷf�Y����ܼD���Q �yGi1�e�R�������a{���HfX2=�}z#����]"ڂyz	����� /��)�K�6�W?��&�c��۸�b�ȣ�5�k�\2��*n�2���0��G�i�_�$�#��>�`�j������5�a��&��N����V��&�������*�dMòQ1'UF�S�����L�Ad�X��1C(#�9�N(�1}9����w��z�j�`0	!F���w5ΰ\�ͱ7�Yr�[�lV4
5i[pSM����d2�Q��{��?�]p�X�3ھ�����ܝ�L�󕔬NON'�>�I���!5;'���w��n׌ɽ9WϘ�1+�#�y�z6=�q��ѻ�1��Q�(ψ�*���'�!	������J�����,�'1���'�(w`<�f���Zk嵎2̴�]�U�޹���XkNm�Bι] ��%���M�>�|>�w��kV�J[�[)g�I�ל�&�ym�����6�y/Y}��jGܝ��L ���p���c���*0���3&8W�j�?H�W˒�kV!d3@
��m��������i~���2�[����(�M�l��{���/7)*l�L��{ͅG���0kS���`�h����Z���L㠠��>�κ%��󖙢�]ì�.��Dj_�#?6+�=wVJuE��Xk��q���Y2��F�"~�� �j�W�-π~=��R��Z�C>��I�;�k���\�>K���� &��f]^��`|.��|�.m�)l�@���7O�@���
Ӊ}.�}K"�u 3�\�!�>��ZO��tF)���)�����߱�]�B������ַ7��x�=�e)��.hr��
G����rs�߈9��jG��Q7_$?��De6�`��"��77�p<Zxπ�{6i���H^���ږ!������Wl��QO�ן?(4:_����.z|��2`�?9n$�� �V�jŻ��}�������Ȝ�u�k}O#F��7���z�T����]?�����ȧӫ��Y#�?rlM�:��(v/����Ϭ���;��\+ �k�^�G��"����ϥ��vFc�"5�η�s���G*��l�a5��[�J��~�xGJ��+-^����G�(Efతo!�z�
�,�x��z����X�|��/����A����$߂����g�n�b4HVrsB������r��r��Z�iY�W�s~�i=���ܓ�b����)�@���#��bz��c��4�[�[���:�lk���~��a�8��#�R���{� ���1�C�4 ��wK!8���KReTkʢA��d�e�#���?�?V�8�y����˦]]>T�����x�z���wf����Yk��t[
Kӯ�b�h�43$=Ź����G,<����H�������!F����83˷�"�"BD�Y���Tf�������JH� d�O�F��un���z����L�_  ��R��$��S2�'nʚ�� �✫�0�n�GLkW��0�5�[�@�j�\��\z#�l�`mz��=b-����Ϟl3�7{�+g﯂�')A�fO䱕�;��(Z}�wR>�2�[~n��\�Ωª��m�'L����}�Y�������5���K9>z	,�`�@����uT�ii��1�=�|%�B��s�d��J�(����Ih����xF��I3��7���+��X�V"��B�r��*�t��K��U�w�L�p
"�+p�
�Z�a��Wȷ��
@�0ײ�)RlH����!'��! �e�a�Ol.O�tw|]fa|��n��kq�ؚx��� <m�����M<�{�	�%&��x������J?[f�Q��i~��ٽ�(�8à��ϵ�(�xeMv ?�u]s�N�ߴ�#� ����LK�i���p�fW�1���ϙ��aP�Ω�B{?��{4��7�e?�H����N�}j�m��&������� �)%�Tjι>R4*9�թ�vDN�Z�H�R�w�ő��:�y��Дn���Loi���ڴۑ���rJ���? �b'E?m;�b��D��ň&m�ʿ��n�@��������dv�髤����kn	 rN�T���-9�eL)g����d��Hb�"���9WrR�� �V��6gL	��
��E�5�L���=� ;Io�����3���w�>��e>ӚB�y��eJ��N�.�V�-�iS�����&��گ�
�8i��z��C`e�lr��6��߫��Q+-W3� ���m���%"\.��hs?�w鵯Y^-`����5�z�Y�F��8��c%��F��5O�g�[7�Y��~�����#g����,��X3�|f]%�m TsA�q�8��A�˴�O)gZIA�/}�i"#E�z�V\@��V��/˶�a�W�uEcEM��֏BTP�6�ȟ!mA?�%d�H�R>2��-c�_��]PՊ�</h?Qx�$D �)<W�a�x^ 2����s�=�U�C��di���hї�v�vA��63U������Im>*V�32cv<��|Td�z��l�=�n�6,�
�׿fJ���q�5�ʨv�<6 ��-�|$���륔��ݲ�L�ͳ a�R����?�3�}�L��<���z�yv�4�<W��a��֌�ٹz����O�{Ʋ`�����r1�f�!���_i*�T��,u�u@[����,1M� �nKU����r*���/��`���Afry��_gb*�2��E��I���`��O�Ӧ$/�kV���$�wL�"��-��t���y�X <7�#�B*�b�l��Ej���Xk�1"� �1��������R�H�﷾$	]��<�H3)�*Ϝ�k�`f���ٶϘ�{�ߣ��g�?���an$ym
rn���ۧ�8�ϡ&W�aHL*�D���u���͈�H�\je� rპ��4k�b|�ج��j����gS�~�JjŠ7���7������/EѲ�f޳fѾJ�C�=�Ƃ1A4��R��������=���V0���[�K��P� y�Z)DD�����\%?ӲF�o]�m��xu�,ٺz�^�����{�ly)���n��W�^/�K�ID%ğ�(�6ݔ"b �k�p�Z�5 �a7��ۭ��țǲ�#�G����1�"	Q�$]�U�ᲕMr�����k���V�	�w�\���fj�dvQ=�R������b�p�rT�r]��,z�\��u�x88D9�7
��mh�D�+�쨿1�K�	}f�Hr�zG�k
h�@�T�|T
�9'�~����=��pdz6�O	�Tg���t�ٲ&�wpF63�ʤ��-�s�|g��Y��w~�	�����o�4� ���x�כ�vjY�f[�p�n�� 8Bp	!����Z)3�"R\�p	�<��#3��9d���r���o?~��������5�/dH+>>~!���P���_b-*���i ����2�c�HEC��o�smd�l��5�D�/ǔk;+[�тg��4�0��J��\l7E>:�+'�L�M^�l��r���6�Z��c�~?:O_��'}�G�v]$�6��R�t"b%X�4e����M�%|��6:/'�S��k�H[iqzc��C��ha��X�̐X��O������&�<�1���Z
3�T,�&�6*�;=}��k)E�sf�b1��hjfR�4���6�ZcXl��A����P�(��]g$�Om�o�s�Z�A.59�wm��a)Uzʹ���~{{+�ۀ!Ĉ��\.���{k���3�&4֏,�KӶnK���s�����V�Zp��!�!��H G�ā$Dw��� �(JL�C�G�>�T����=",����fp��2�0?�Il�����w���./��_�ɃM��˒L��zʰ��B�NY0	�<)�����t�M�?���ݍͤa��2�[�nK���4iZ��X ��Z�T��W���2��#��g��G�w�<~VbJ��d�y)��C�HX�j�������(1��^�!+����#���w*�'�D�vz�Q+1=����V�	�^��e֝�&�W(����)֞�<o�[��J����=����؟"[���n��y{֙�-9�EξRBr�3c�" ���C�+�D�K��v�+gԉ�C��&���;�;�%�/9������'���h�8j}F-�d4Q�yێ��q�H�{�FH������QWK���<��kf��v�I~�	�l���k��F�ˍ\���f!Kߎ"�{9Sk�*!���a8�&S���ض��fl�v���l��0��̷Ņu�-g�P���x�Zb�#K�e���H�@���!��#���w=�
�R��z2����; 4A��2����d�K�Z�������-]�M`���� ۻ�?��g9�JLH��L>��P�QB��S�g��4�AX��X*k��K�P���'��ǎ��?� fӺ���1,y����_D�s'�hۊ~�h`�z��9 ���Z��/����[�F8֢j��z��,áٮg�a�io�����r�HN�}/�;#��7�=3�&Ѹ�ֺ���A�1�G��0<�����)�������\�� Q��{�<�����R	�0��ZҏE�n<ϖG��O-��Gs��#m�? �up�^x.d��*��`90х\0&�ĕ�[����@��N`����=�v�~����y��p���ccJj��3�V�P�)�M�N,�aS(�OQr�x,���k�pצ� ��,���l:BV
���ɥ�pf`�V, �f�3Iןe��l��|m�����d��h����/8�(������?�<ohޘ�fL����=���w.�S� bi���m��)�}�N���ڱ���'��2�9����hlʾ����z�`���=�(��N�T�0�������ѭ�a���j�٢����oy�X|A��os�+��HQ�b��%�;��kFtź^��Y�^�X�1F��r4xڢ�o�[�cs����; Gށ���W,�1&�k��,��m+�2�,`�0���g�um����
��*F�7��Z�8Ѯ+�~X���Y���D��c ��Y���2/޻��"������E/����|��M����ϯ3=��� U�u,Z���d0g|%������j9'��a1v�m�=�RD�~|��>��O� <@ÿ���2O��T����O�������K�u}tk�_.���%����nM��ܑ%��=!M�=5�d�F�z�?"�
�}�|E�$�O���+I�3��~X�o�B�% �BBQ�=7����{}�%�" *{]�Hב�)r9�����ϒo2e�>0�\m�<� �����c�uͭ�pc�s.�B/�׮
T�M�Q���۳A��XH���$z�B�&���v#�tF8YxQ�5���ϲ�)��%-&#��ؐlS
a_EE/���3�P�p�Xr�r�ʙ��#�6yo�����O��J�#��g�b>�\���QJ$�l-��=��Q��P���ea��s�ҭ��@��U�7"ʻ%j��j��Y*�^��z�!m���/%e����(��'�����M?S�3��֘Yʊ���k���kAF�ؾ���cQ���Wȷ ��PJ
�Ϩ_>�MS�-�]|��7EHC�,�9+M�/��Y�(G���E�b1�z�ҠV��-�1��J�-���#�K���>ϜoUџ���7�Qt��X��{���R�����c�H�mf��B��9�n�l�Mn�ٷ��3��2=�à���NxN2�^���H�A̯��r��YƱg��J��5��\��s�_��{�F�	�ʭY����[��vʮ'��r���ઢ��)Q�5ʜ���.=?��\��slQ-7�0�zϫ�#�@�D��%�	yo��^��FK�Xo���rYp].�,�˲m����n��dD*�/��ŗ�#��+W�H��.�%�_׀�EaX��~q(Q5�bL�i�Ӎм�c:�pK�\� $r�����l�S!�M����Ѻ���ƑX�;����լe��'�4�@Dw� )�v!�聆H����(ʿG�=I�{�|j�)�����`��y.�38"вǣ������1W�#n:i��E�s`+��g�\����\:�k�w�btf����+�@��"�=�l��z���^˒��O����h�z�e4��q%ЖE�/�7�Ί샴 p�!Ɲﴕ���vN���ww�'ڑ.��-��+Zһ/���2��  LD�C��r���m������$x�fn�M��sz�m��Ϲ�s.����_���w�V�a��;�˘L��y 5�$���b~���[À�k��8���6sYX����"ҷ�M3|��L������܇�k���7+z��g�1@��?[v �����;S����6��;�|�ane�o�z�<m��`��WF`�edb��]���e95jE�N0�Y�錌@�u���=�}����rͮ��� 'd���U��0�����p�u���#Ṧ�%,�ZӣE������R�G<��͉�����s�� [}��#�0��g;{vNM���sb28��� hW$��Z�@3?�r\�º��ϟ�����:�Y} �Z��l���\5����%�F�� <�O��JuP:j@f���F��
@�3G�4�H����5�>c�]bm��g���.�W��|N�ۃȫi��<��g��IiK����mF���1ڣj?��V���6�&@�h������ʈ��߱����5�8��@�h3�A��FW��L��g��=:���?�D=��Z�����MCd�C�Թv�'0�gs@��1HؒQ���sQ��Z����JV�&OB�'q�ul�}�q>���� �ϖ2��;x'�=(����s�Ƶ����c؟�Q���y��ǲ�$�h�{�壢5���d��6�!	`���5�{�M��ţgGk���}��5Y��I��U��f��Ŕҋ	�f�EQ+`�ܔ�]e?R�fX�#Ӡ��f�f��[��ϕR[�r��Gǖ4��>Xl�\W��) $�k�S��BV���������#������~��2qx��t}R2It��:�R|��U.w��T�����	&�/�
>α?�0�s#K���d���d������~��GH����)	�����7ep��bNLer����aL�HX�Km�r� �� C��_,�Kɉ�J]�X��eY�H�@mk���*�(��L���w�%��Z���h�l��iN�VKz���1��s��?����K桓���g�ϳ2����f,�>G��V+�j6����^��#�;��Ќ5�[�I�c%���T��(�������S�my�3D9��j�^���'���v�}@�_�i��j��J�����ëWk���pދ[A[~�|Х�4����,x��G,�uo�A���FǤ�,C�,KU�����l*/A<`*�<���s�&;����}D�߰跓�1��<�=ХVSȭ8�T�X9��C~�?��[.Ŵ��E�.�PC�~J���;{��j�� �ϔj�P����>Ӿ^��5����k���[H��`�Ur�,��v��Rl�x�O���p�,`8�jɳ����G�f�����<͸��X��]cw=�`ZJ�ѻ����{�yy���z�4��vS���]�89F��1�ʕ�ϳ����7b��u��5��S_c$r����g��΃�<O�=n�<y/G�1&��f6��̗$��_$� � �LO���J֗�@�%��tX����	!֒M"�1����A��Y��L�������ko$:Ik�Y�Ѹ�&�ܳ9?s�U�`���h8j�H��$�#�@�����<_��M^Ӫ�(�cfc�gǥ[��1�g�rx�h�>zV=�zVxH�y�0��7=ӯ���`"�^Գ@��+3��Hّׯ�r�K�S����:M��h#}r���M�XM銕A��e#<ƣ1c�\�0dLY�a��d2�tD 9D�C>��[�X	�Tpǖ��y_��^��"�钃��K�d&{^�6���[������@
 'V�˜)?D|||T��z��z���L)%Gfl�7S��+� A+�%G�?[����Z��ƫ����W�"��bgDc�~�h���e`K��
&3{��D[�/�K'�Z}=`.e �	���U�RpdJ����E���P�,'*�8l�9c�9�+�=9����
��gڸ�"O��Jyz���l���c�������S�Zn��t5��Ѯ0�d`�^�@���س��G��I�;��{$@���%��S,����f�@��^Il6/d '�D�S� �˷�&	��]�1�X&G59{����b��"�<J��ǈ�)f [�v�DդUϏ�&���.oW�Ń��q�3!�5�W�m_��O�B�1�"���D�+nm�������#��i��Fo1H��nd֎����Y-'�=f�>\�L~�p�Ȧc!�|!�0�������~�H��"�̝<�����b9��C�b-�q`=��&$�yNO�
��7��
n}����g������뼏,=�N�?�h1Y3��4fi1gY��Z�����=�9����c�� ����aS��+Io���s#ztͼECB�5S�>�T��1%&3�|+g�>�Fi[�֚�]�<,8#��(@9R�	)!9jbIʗ����el�b-%΢�cJ�}���\�}6�G����̌�0��gh�y��rn>4�u����oS�E�s}�b�	R��3݉��i�~�2�����Z�YU��%#�^d�DX)�$K����Q�lbՎ;ח�K�yϽsG��ڰD*,ܖC������4�S��j��PJ`r�����,�+VNQ��3��%g@�y���U7)��J/Z�l�s��#e���Y��6���4��~r�=%���^�E�ߒ
�Ϋ�l9��h�* ��Һ�@ӕW8"Dl�=p������=��f?+y�¸���&��'Dʿ��B���S�1U����z�1��Bn0��#�
�����*{��^0�Ģ"�P��r�R��L~C������}g�1[:b���Q��p�?��5�Y@h4�f|��)"�����y=.��x�������߇fqe;3�`Āͼ�G}:�J8+�Ys�n\�P��q��Ļ���(�@/3��&g�g�X��ր� {�;����3]k�ۗ>�y:� r�Bf9*~�@��o@�s_f7�H��d�5�bϠ��������3/�.� @��0�QG�= �F���ll�kLS}P��e?L�V�]���I���(��ޔa�;2�l�h��6>��#&�34�Y9��~��6�]��&ɹ�V�gIm	^��d��\�D�=!�(k�1���`��M�].H)59?%0��E�S��;V*�< ��{��4L�`Q�~$�a<�߃
qh�����#�g��߽�Ao�7˭����3k_J�<s��B4O00�Jf�Q~�|�#Ʒ�����۰���?9�zm�ބ&�Q�+�?��,����?A>��ż�ErH���|+<2�쉶��Ω�)���<bHp�0�H�Y( �7�
�?���i
���	�ݠ�Z��
B[�����zcך�^��ސb�y����2�	[��������e������}�ۯ?���ˌ�M4
@�����s*�\E�W�ot�Џ����U��yF��l�׏�w¬�c����b9h�F矼��1�=f����1��k��ɡ�
险{B��+ί�C�єg���>�.hf�l�g(�G��f&�c�:"������o�]<�g%��Cr�ע��)�w|�����p?�}��/��e���^�Ɍ�������)��@��'=|�* ���!0�JWy@ɘY�#�=HS�������?��;�����Ͽ���_ ��}3;����rԄ��0hJ���;����9 8x����%�4�A�F���js��ҩ�'�AZ��C�ݚI^'��ɎS�v��!dU��[�k���#����lm�[�+M��{xj�E7cB���a+G��g�R���J�'wy��W�c����}�{�������<D���Xϴ���wt�n���}䓹{�'}"5�㼧�=��e�G+�P����u��qyf��_�����[��d=����V\XB��,�� R��ON�ą]�$��R�� ��~�l:�Q���G��7)D�ir�+�% �_����o�\(�Sʑ��6�9�[<8��V�jdE$��jev�q�y�$1d�k2����^�bw���ծ�k���  M�V ��v����Y�-@qo[������&V��M�Q�������'/vm�"fj�B!e������Yc[u���U�\�����̳@��GL�Q;�n���>��2b<ynܝ+�`��Zm�;Ύ|�geg�a��� ��O��J	!�:3ߟ{�M�Z�\�[�L�9p�ae۹��{�""���Gu=��f&ʀ�9T�6+��-H��nJ���$��D�;'�4��O^c.�O����zş�\�>.�6�d�z�٥� �f[�i�8l���Y�3SF�ە���yH�%Q���H`Q�a�*I5�w��q�Ao-��ybS���Y}{&���|��|���L6L6K0� hA�L�-�l����-�7�O�*��Q;��� P�io���3�#ڏ���:��0R��(Yϐ(���o8�T��5֞1��5x�,Xi�>Kz}����:V��=Y�f���a����K��S�i�K�����Ss=����7e����R�߱W|%�p���s��a���d��?Y��]���܀I~��d��+���.��������ȋn��qW��.m%KBN �#9��y��q<�D�M`+ӯ�"����p��s��k5�8j3�NY����B���Z�{@֪Mޛlr�%����L2#,@L���Œ����7�m�Cd-�# +j�U������`v�bʇL�r�����.EW�b_D-�_��ޒR�)"#��L�k�Jb�C1	:��y^<�����<�z��8�6u�!�~v�ƴfW�wV�%"j�����z��3�ן����\.�K�<�zF���g�a��T�z?�����z��[V�
�G��������뷴x��V�>�R��%Ou.���SL ߒ##	!* �%1��\V�F)ܼ�#�j��1vź��"���p�\r����r���������e�q����f1s��`y�	5&�/����'�ն��D�Yy������ϟHnH��iެ5�����e�yJ��B��!w�lڙ��Z,_K�����A؏�^�e�3�����hS}֫�"E���r��L����5��y�����tѐ/Srm�4����V��t���ɹ�Mc� �E���0hf|3��.p�p��[�(���s�7G �H��Ϥ�Ե��Q��ٔUR�bdU��ϡ���,f2<[f����,K���@,[

�޼�����L����%��o���b$MF��{W3^�"y.=T<�'w׏�fj9f}/�x��*L"b����T"����� f1	_;���% ���?C���r1K�1R��S2�I��T!q����b �q��bZIطz���3�]�R�<?ÌX���w��ڒ�c������`v�噛ٳ5�� �����{��L9�2uO{@�]��f$Gng���6##@q4�z�j���%x83�Tz�fo�qlBa�׮�?V�o5����L��Q�gm9�z�Z�e�k�?�o% Gk�p��&V,�)��]�F僩�ɲ�5���`��w�6�u�m��ϻE3>A҉�sφ1	H����'P�_T�!�Q����Yd}�U��Ã��Y�6�sJL���y���;����5�z&���=�:_�?ƛOȔb�)��Z�Y�hʅ�7J��z��nh�3U�>��|��g$AV��5�ԅo˽ S2�H��6_%��;���x�
�n��5*/���m�im�:�d
��ϕ��3,��D���K�9�ƺ��i�y�<�,ɺƝ���GpK��1�g�@D5k��q����S��Eo���(-w2���ϛ	*��;�gvW��YǬk	�<��;$�0S��lf���R�`�~��,΀���E��J^SV���/�B�X�')�V���}BBL��R�k��"{�/��f�W\���y��J�~��������K1�j��p��E��ք��i��])�6I�#�ϭ�sh�i�V*p��U���̺�&#ϕmXmk {V��M�9#���^�/�=`����ce�(�{MR�����z3�ƟfN��ܛ������ؽ7��e&\꾌�gM���G�<`�h)���]>��pcf�-n���=l����f͟W3�=��N�o������7�������2�,+m?�{�1X�l�
�-u(MK�3_#2���y������]�6��^�2� ��g�{�Au��@.U�9����SdI�Q�u�ȝ��
y	ȼ�>�?���kJ; yV,s����
_��X�w��;_�Hr
�=�_陾�z'd����'�2��wu���D.�=F��NX�ߝ�[�3Zhy���L&�e�d[��ɦ�$�>>3���_O���b�dµ�"E��Y&ǥt,=_5��hKΘ׽R6%X���}�LNg��Ǳ��nD�9iv�r���1��
�[?��J�d��&����rm���ς�@k.�D��J������G{�&_�넚nh���H���4L�
Q�e�0��hc2s�
��K�EJ�<����f����% 3�\��#%� ������S�wF2��	S�D%��׼�d�]�D���γ}�E���M���KJ%�Z�OƈP<b(9��H#�H@�kK`a݃n�Ԣ�I��Q��f9-����2{l�p_!�?#s�X�#�`ȑ��k`:��<2~zs�b{2�*��j��"�5���� h-%��& R���Z�}e�e�Ӽcݔ�ɫM�#�|�����:�˚L��?�/U�(������~��sE�d�oc?�)��8��,޻�;SZuYG�xari�$��3��VRj�宀ˍd�ʘn-}/y	�$��$sI��,M��g �f��q]AރR� ��b�wio�׷�x,��>����t)! 6��PU״!k!c�<���b�3/�L:Gm�s��:G}=�N~���IV�aVr�͑�^,p��ĉJ�;�۴�����W>Sm.=#[*�3$M9L�:��^@K4�k8Ú7�)�aƏ�jWZNzsC*��u�媵�o$���}3&%�$",%�������A�/�2?�F2�̼B,�\~7�$��'������wx��P9���B��ӿ��4�驌���;�E���@�:�6sw��}���7�x�O�t����"_!�Ia��w���?#E������h#���M��,�9�<�R���a!�Am����~Y��G�a�PSs)k`��ǘ�9Wq0�f�ф��[f�ė�64=��m[)��fzd�}��T��q��"/Ɉ�6�#P����m��ĭ��&�3U���k>�����h�ɭ���`V�.��)諭�A�R��<�1�Z�:�T*ֳ�JVe�(a��tҵE�	��\� �6Ǘ>Y�"Gs���n��~,��X��HI��"�{�?"2���s�G���=+9�p��：�g(�>d�^}�����i�m�1i�e$3��z���3zJ�H����F��ъJ��^[͜����fd��"�N�d,B�L�d݊8��>�w��l��ᢏ�,�Y*�Kp��)6���@	*ș��Ϭ��g)�쮓�� �T�i>�����5>���Ê��j�P�E��\yAg���$��ϔm�k��)0Z-ĳ�o��68��a�&���@�ha�W��[�s$G}�Y<���*��+(����RU�d42����J��c����k��x[Bh͒� \`H~f��>��X��gS��k��3��Ϭ��S^$��$=>yLiSvo?2��U�β���պ3�ό�>{��\����_ݬ&u= ���Ǜ�h�S/�mߎ�`U����z?[��"@�ީ�l$e���i�%�����̀���Y>>>p��k�� �x�3;3�􋱴�<����!yJ�-��N��Ȥ�M:�A�e�Z-R[��>	$zb%�����3��#�����0E�\��펗�>)�d?+�sG�gsn���@3�� y���	�#��<�&f����v���gm�D��]��a���+�I�ji�O��#9:F���+=uƴ���eOY=r��}��}�5��^iT�oy�]G�]N}d�iXm�Ȃ��q�Q9W�"�L��U>�,h������u���`�w�)곫���"2�,�y���Y�u�m��kbD�!��Xl�f(?d���l[�����Er��U�豭�X�դ���y�#,�#%�=���:R�����b�������}�������̼���LR�5z �l� bb�bŵŹ��/㙴�g��#�ɣ�1M;K(�}>*)%��[�������9 ��e�X ��r�6BC!��~�Oy�?�������kũg�>ۦ<��|9�g+�+sl�)���qg풄	��$�|-9	�}ƪa.�e��|�>[�d���-����*�6��lg>���� %��9�8g4N��4@�w�����[����&�/�;dހbB�)����|{{��?Df)�<��t�\v�3&�%U�ܱy� ��k���&��Z�f.m��η��)�8�b ��d{`S~vh�4|� �~��w����=���@�3݆lg�䱊}���}���Pe���o
���u~o�����r\�39���Ҩ�w��1\g�ί�V�B�v`y6�d)jg��5����W�) z^[`N�E���۳Y����S~F�#�'r�ւ�O1�zNs�ˣ�������$I7���ZtII��d+5���#�["F��ҊBT֤�o�2�2�I)�S�#�3�$b�R�]"ݽ�rP����y�<���y�B1s�F�$|�iQM]?U�d��9;kH�Ӓɟe$�ND[�����d��HǱ��G7:k��@³�g]ۺ/�8��Ѧ3�]�DT�Qxk��I��Q� Ԓ�����)�j�����̲z���p�1���C_�"F̖Շv��9�Zʻ�~��Hy�>�U,��R�1 �N�s}�,��K� �bg��1��z��?�s�@�cb�$*�%��4�v������CMY�@S�5}yQ
#W4�}��� ~�s����9��A{�����e-�����ɡ� ��5#D R�c����
k�r�iVƒm�ҎI��L^����>�=���Y�1����UZ�HtpV�n���gs�wl>��Y��$
 �T\ߣ�M��&���3���~>�2���HD�vo]_ʈ�����h����l�#���ˌB�dҿ���=�&�])֎bU߿�aU������[�t��3#=�nSZ f������~2IęP����lk��U����M1�y4eNKY�R$�0�j��\m(��g!���[�����'SG�b�kY"�m�PQM=���Q.2��4�2,�|�����np�O��< #�����Iאb���S%��	�,�����3p{f����̯I��L�caKp; �;���r�H��注[6��1��Ly�^�wbHA����`�U@����#�=#=@��#>�����u�=�9�כ�γ���}�*9Z����{��KKIk�7Ϋ���#gޭ�7�}C�3��6�[S�5o-?K�X]� ¥�,'_�n���u[�_���8R�u̹�$��^��3�T�>�O��If1}-l��% s�E���zE)�3f9��±vR�4}����å��B�M@���)%���'����x�>�rr3�]�\�lY���K�3N�q�<�e�0�O�`�8
]��:2)�zl�,8!�Z���u]sT��/K��Q�`a�؞d0<f'SJ��� `Y�����u�fzO�s�!���ȹ5pPM�0�o俦�o>������}f|���h��m�*xI�-Y���AN�F/�c�eUHmq�����}�z�����Y�>z �|�r6��,@�w����P����,�<�zL������ݩ���1�<��<��s��}��ǩ>~�|ٗQ�.�}]�\�٬O�uH�Q�n����P�o@!d���� �q���e���3U^~-�������Q!ΊOf��R^2S
Xװ9X��P��"�f�Y��oo�}�imb�.�4��rA���k��>r��"��J�.g��^��b��.۲L<�$���G.��ټ{$H��P����wV$#9+:O���Rj�Z刔L}���d����]�f�Y
��0�����=K���}s��TS�P:3�v�e2�3�����rt�޼=�NoߑkxÞv��|uʢY���e�)�7)e�T޿c�1�]�Ւ�&�RVkkjL� ��=�e��z�o������^y��(?trmI�*��a��ixεţ���~P�KigJ���
&ͤii��a����:���v4ȴ~>�Q:2{Y�٘�;�Ç���Y1Y�o�8����\7i����#����kγ6��c�n��� ����YkݑX{нJĈ��vϐ,����G,XA����DQ2����Z<�*[-�;�d��v�m�ePY�=ժ?D ���1��Ώ���튷��j%�N���*�ID�/��z6s�K��$���U�z��3��b�� �}6y#���Xܳ��] 58+�TK�is.pl"�
�A�!2�r�,�,���g��m�
E5a;0L4�g�}�����P[Jő��l_y�!�"KV0�,I՞�e1-po<���{E�����z-��%���#�s��8�gpvK�b}_׀��![iS����������v*�d��$s�"WbI��&����b.�%�m�����Нw[`I�xc�^r	����ܴ8����y	�yβx,�_؄_Cr�o�����O
�YŞ̂Q����*D:�|P���,�%��{L�����Bwf!�I��aooo՗4��D8��h_��X���Y< S|t�2E��b熵�嵀~nD�X�>��&r����Y��1�i�L�=e������v���,&\�.V?g��9��f���&~������>2��Ɨ>��A�j�ʓ)O1V�I�����?4�6*z������z}����[b����XB�H%*Y h�Y��X�,�s�=k?1Ȓ=�����q��� ��yO4�_
��x��#�R�)MP�s�rJ�C��[y�DsG������].\�����oW�$��JyM
#G3�U~HM���`*��% 6���6L��S�H"e��.F/N�E�^�l��X��#R��E���\�����f�<ۤ$A�Ws&�T�َ���1$�f�����clXFK��g��H�]E�2�.*���f���FR�\F�%�Z����=ŋRJ�,h#��N�B&��뇔{ַ� 2c�� �J��M���~P�H�����#c���VR���k����!�_%|-ΐ���Vs�8�����$�\�
��&� ���ٖ��D̈́缘�Z��#�䑍�̹)%$Q�q�_t�����=����дdD��k��^�3�c��d��ޔ]C�D}���:��3ǟi_Wa:۞VH������\~g��ѱ3���<G�=�bώAΗ\�J��1D9�B��|�,g�5 M,��b��׾�y�QT�peJ �Q-�rJ~�9�<��w��d:Py@3����"����z����R��0�K�����@�qլQ�!Y>���++ڛ}^G�hO[>[_���leMsS�+�F#��d?H���M�X��*�7ir�c�2���ަ8�`����bѸ����
,��ƿ���Ng�E�Y�K��
㶉����\���߯G�"L�c�Z�g?��3���v���w�%+H��D�_�#L�)f���ߌQ_�����cf�#DG���$P$ �Ƴ"�6A�%����'�Ny�_tn�/[Lb3kJ�!���'����)d�����|o6�:�AlF��=�i��<ovw�)f��:�-�O�t��cS�e��S ob�
;"�e�#�Z4gZ�&�\ÆZy�k�$˖�0����,���%RY>��F>i|�%5�k睎J_r#�=}:W �_s*Ӽ6�YJ���S,��jc�3�P�\�~eK˳���*yq�?�L�Eʌu��ʹyd�� �ȇ�E��g�R���k��@T�'�����o�_�������Q�ޣ��?\�GZ^��h\)G#���N���-��=D�7#?g�_�#��}/��֧�����Gx̊6�$���8����d̓���!�����~m�� m�%����L5��s#�Ե��R^2A���;$�!�|Tb���a�4끙uc3Cc�M���nOW(؁<� �f���Q.�c�#����:���b�k{��~�4�ؒ���v�3���pp�{LY�Y���q�ZcO&�'��*=#�q{�z͆�Z��d�-&�9��Wp��#��w� ����D�*]9+Z:�#���Pa���\b@������G��k�M�/]��a���끃����5��ψ,\�J?���G�Yt�$�s�u��K�
'�gV�� ��p$� "8��/�e��r��z����.u�w��E�;�j�y�o>3BD �ۉEMU�}D5�J)!� �<bpn�~(kXA�k��Gq��[ ��>�x弗�"
c�@���0fe>C�9�-ϛ�4����	v�nv���=���ײ��
#���J,<&���5�И�c���dcF�5�.=y~��o��G����� c2 �9o��Е,�rOB	�48��g)�G�fל{|���V6�?|�d��@߽B����m9VCaK���J�����`�H,��n<���'=׀g��z��,�yfI�uD$��UFQ�/k���c3���^�0D(i�Rژ�ܫ�5K�"��/��?~�������_�o��QV@6k_�01t���r6�MJ�k�J�AJ��5�ݹ,ٺ]�w�Qh<�e�u�I��&�n�ZN��MB��3>�_({}�1��Mv�GK��7���@�0=#���PS���'f�b���6~5�_��]۝g֫�,�����Ҵ���b��Y�`�����ٺc-'kݫdc�3��h �a��{�=�ta�sߪ�tF�ԕ�f��5,��ࡤ��Ν� prq
�����3�����(�Iȟ���v���%��b�n��i�S�T^����ǽ='�(f�v�Ĉ������_�#�I~V>w��-.�׷7�������������}�DyQYɄ6���dt��t�=���سm�n+-Y�]��������jE���;D�/X�\�Ә4���$�{d3YQ�CW����##L3�)�@�.�}�,�	��ͦo�~�1Ҳ_bQ����͙�����fڱL~���d1��˔�Q��<�������w�gJ����A��g���Tn�V=��2���<��B�@���7{.���н�r�3,�L���9+���5Cj����r�
���r�>�݇P��'�q�/.��l��������ݺ��4߫
u �{������������4�Kj��g��:�e��_�)E�SŲ��<쐙)U ��/#@�0���hS���X���r�`�\qY�������_F~�DFl�3���  �����cD�f�zjw��7�����1�TEgDG��0���m[�o��Ų�sgA�hT�9�?�lqoѷ�k�z�g�dG�i�ŏ�w����v�[��]���q)�$� ���dG�f��RV�{`]�r�+0�0�������eF�)$�H_S�ȧ+A�=&�g���+n��~�3�Y�q^�t��3R���M�=�f��c�T?�{ݷvd���}i���x�1����kXB��{�9 	1d�������qIaGA[� ��o�w�׀�C>!�'O�qHwڜ�P�_�d'�vt���x�$�'��m�|D�ц��<�ãL����?�Z�8ˤ�?�3�7r�2ѓ^
��1i26��A�f ϊGG��"A�L_�=f�!ҭ`T�]�iǩdR�ְ�y�Be�ke�Y�V���`Z	�����j��Yz�p��g,w�~�XН	|�z_I8l}%A��[��_�L�6Rݒ��Qe�c�!"ƀǾt$f�JW~��u@�\��K��F�\�K�;�8N�t���
yMş�n/*����~���p)]#z2�)�,��[��l߭ϳ̵�c"����a*��3�z9�԰%��-��n�b ��w�1b�$�c��SR�Y䏘V)5E�O�K2SŦ����x���MX��3 $�X7C"²,Od3fF��d�k{*��?�9�L�G���1%x�$q_w$����`�m&��p��Q���)" ��\�����3�Y��2�����ao"�Y��^S���%k��8'�RX}і.���q��wM��j����,,���y�~Ks4^�fָP�{���u��t�1ePYXNJ��F��t�%���_�����q�,X��% �z�fPy[q���'"ĸ��3�	DM�ۿ��S]3k&���*)%�5��퓫�y,��\.K����P�8�����B��M�M+�>~�y-�� R�A�-h��� Nˠ�##x���w�#���?�z�6���Z֤�_��Ϯ2��&o��ˎ&&ȟ�AB܆~V;�J"��O�)�-��}]�f8b����
��;�PN%}�XL�r4d����g�&a�K�f]z�Z|�3&KNX�b�s� �\�)5:c�����$+�s!�nG~>�]��G)��!0���Af�Xi��\�y?32��Z�]���J	�Y���6ꯟ:}�n���c���ϳ��S��sF���f�ǰ��@�`�n���	�`S��z/���y�@^�Y����M���e��9�a�L�p)-���p��sG1�����~��5����ט�)fG���r�b�E9�����T��$B�-���5�-��s-X�Ǘ���;*��&?��N=���l�Z��0�߯��õ��k-��q#�4��T���T7Z�?o$=�"���Έܶ	�&��L����4rc��Q�")2�o�g���LV����տ��ʍ ���S1�k� �'=�{�Z��v�؈-@phyV�3=��<ػ}~�;=R�/�Ƚ�����g@�T�z����,��[��\x�j���n��~�?�\BJ���Ny�ݽ�ԦD��#&3ƈuMP3��F"D��D��ti-&u��{�,A���{���J!���|��,Of$ p�\���s��O�	E1it�* �W4���N����N�T�J%a?Z����3�[�sꍯ�c�f
c��l�,�8�3���1#���"��~f�����}	a�Jh�(J3�l��M�O3�Ԣ:#�BTNYh�Eotl"�J�c5��:�?�}��(�hc9����SI��c�ˡI� &@ٿu����6[�D3��2��x�0Z@N���§��Y����ޫ4��@�����זo��u��=K��g+�[�Xi/�s�΢�{����$"\�W\.8��I��r���GY|2�����+�CG��)��9,�KU�c��}|��ￛ��Jy�O����m��F�U3��x��^S�g,�_�~���˒y?����h��h`��-���\�0Nڌ��٨s��nE����"��R�DU���m�ь�#�7�u]�Z�o��즾�,����ʹy�w&�f�U�X���l̴Z�CG%�4���"��(z2�� S��W�k4�t�0k!����%%Q����ϝQ��}���ߪ��f�l�������զR����eg�y�z�s��c]S������.�{_��J����B��j�m�F������4�����ϩj@�����{�����.���u��9�r�d&�.��z��r��rŲ¦0�`E�'��[��+�v��E]o��o��eL������ b�����\E�[M��Jvn}|�ֹ,�����y�g�����DY��~��췒�$3��6�2�0ȍL�d�$�X�&��[�t��g5m��@��>z;��ښ�56�J��V�d�y6��J�_$�A���X��یJ�+RvT�X�^�D����pw1BqHe���u�pJ��n�uF��k%C+!��'����d_f��Q�F
���L+A#�l+�k��N��# ��29�{mn�W,fR�ߓ{v�kJ (�l}�\_�Cͱ����<Rpt��8��u��vu�x���=���K��1��u$�h�4��$��t�����?+'�|w�˂�m3�{ﳙ[��׿����w||| ��m͕������6��������w�x�T���gL$+J�y�v5h�d����KyM2v����	�\}[(�`~xQ�<C��"º����م�㤧2����6���۝S���>9�d�Y�=�=��8K&c_����s����J��;o���2�_�\c�$��aM�#�Ms\H�gD��{Ͽ�ޫ9�ຖߕ�`��}�3}�����=��F�
ō�tg����ϧ�����n��H_l)�{dF6�~Ї���4a)%�^R�
4�Zq?+�hp��J)յ][���c�n��'�J}O�����&�yvHə����E�8R��q�������h˖�\��l�f��砦-򥴶/�2'"lϫL����g��mr����U�G^2�w���]D]c��>�
�����Z�Y0�ck꣉�,�����̗#�R�ۤ�"�X�0�4�sX׵jP�u��,����2�2	���_u��XLu�#��E�n�MBr�4>��,�ۤn���A�c�1�g�h>+:�aF*;VXi��Z�9%��|t}aot��5�t��V8d��!=&���#ʩ���GK9H)5f����+�wR��:g$=�r�e�.һ�%��m@�,	���	���h�X�]۬sFl�5{���Ε�f��3����	�A�}F"�?O�U��&�p �s�<�b�Jac�	���u�!
%(b�)X�j�42Z@l,eq������/���P7l&��eG��/�n\.�+��+�ˎ���˲ �P�m�wU?,a
���R�-�쵽������8"�� +/�T���e6c���YMqt��=�뚃���!:�nK���������Q��Ys��{ɔY���}��p!�0n��&w�4��6e����2���H��E���d��{�YS�����UQ����w�{�'|@5S�b��b�����?j��f���a���:ս����#�\$ʙC4h�]G	�b�dxe�Gs R�#��t�*������c�+���]�v��[F�D�T了��UF�U�*9�Ad�c͑	��I&�J�V&�h#�jO�h�=#/�k�����.���	?2{薜���k�X(!`�9�L���vΞԷ�x����ߐR@N��s^����������{����ag~���Z��#��u��^nx�G����HO;����h��v����B�7�Lz����Ё:G�CX�~���bsm����M�5�P6T�ǲ�c=Km���˹%_��I���ٍ���4��?R�dd����k��[r�j�L�_�dye��R��k494U�We3�O�n�{/*���Ѽ�"����{vK��Y��<"���>z}���})%CW��]S�/��h�c���l�{�Y�e)N�v�X)z�Z'�����T<��=��A�������7 �-��}BZ	���������r\�c��k��^[�coY�>�1T�3�T#�[*�6#J�����2ƈ1"G��,�w�F�3
rȐ��	 /@��p�@"`��/��Z�6zL���W��#B!�v�a]W�n+���G�������~�T�S���@kN���c�j���S ��Q��'D��OҟS�c�3#:咔3 ���GbE���Q��f�� �����c��Yjj᪐R�+���ύR�̅�wK��cS�}>Β�rDD���W �D{l�j��D�7�S
+#ֹ5�E\sČ[
�Y�W'S���M�����9�s�d�ki��>fGk�n� h�뤒�cd-����5�V$}No�}NR8W3a{>M�P�{��:��V���<�������އu��Z}AV���HHpp�HΞ��=�R@�R@f)K�}/yMt�w n��?���}z��������H�w+��״r�˨4��6�� o���*pDX����E-���L�feԊ�8��U`���&�S�P�/(�~�a���ג�*�zV�<�^GIw�s��xv�$��mq;:�d�Vf6���˳�V00`���fL���8����  [;$Ӣ�٧:ۏ�G#�{�[�fe���,��v(U��J���S�eG��~ޓʔ;� ��vzJ���7L��m�2c�9��KB��ܫ��	�:�-�A ��ǐ�#	��j�]^D3��\��sd�w)%|C��"�Y6���/��-�����Z���,�#�a2e��V���{���R"�Ǐ%�Lsk���B�#��4�^7�����h�t<9��tn��_MF�d� So�����6Ww_��{�����{�t{���:ꏾ��T.�8�aa��L���&�Z��v� �z�:����dfs����n��g�����m���g=������[���Y�Y?�1C���:�
I���u���{� ʜxp�5L���ѳ�Yr�}��'�w�bw}� >�Ơ@�np�ؖ�M%<bj��u���@4R`�<�=o� m�>�����{�}�M�����<j�}.��E�����r)�z政^.���,��.���`F��"�q�ݰ,��?Z�Y�����\.Oi-虑T�)��s��ϥ�'P}3�7f��9�s�*�&m���CB�1�{L����Q-�O���]j+o�N�ѻ�� '�3�������b����W�{�iv�
|��c��>�����w�X��)'�=𥝑Ѧj���x�\$��~g�l�Nq�]�?�w���LP$��lV v h��� �
���������ZeI/kB}f
�U���3/�h:@�7&-�>������Xc舜1�G(�����<��ϼ�# �&�_%l����K߶�Ӑ����)���}l��!�7x"\.W��$�|�D۾Y���T��rD���R�r��\��-�D���w��D����5xw)�q�(]�Z&�o��B���#�.r�vo�[���A�E\o�1��D�:B�R�>�U�B¾I�'�阹�gC����L��,�I�0H�
Y��L�5�j�gD']�����{�vY��}�v��O��}=��gUn���wɛ�� �#�bVzc��ti���.�^�w������4\��J4���+Ƿ,3	�S�0�yd-�=Wn�2S�����H�x�x���J�?Z�v@�À�0�G}�G�zF����Z��g"yF����; ;NG�[���r��~t=�\.�s[n�H�\���9>Q��t� #"�J�E�gy��,��)>�������eR��9S���D�5� O�pԦ+)}���]�3�sd����^�%-μ#��^oT�LbG�Fk�G%l���A�Y���\I�?[v�פ9{Vvm0��8`�W����t6�Qt�2�RX1i�>O�P��S���{.��zp4&�@O�q�/�ܘ�U.V}}�ͮ;�+Fo�
�l~X�d�#
L2�(�̰�e�R����3	Ѻ�X֞2�SJ$z��]��7�, ��w�z@"��2v/s����9�P޳��<ɌR(S���, �#�	ٲ����fyS�^]�'/�]�p��L�ͫ9��d+S��R�5�$X̦� "@m޾��H��`��3��N�����o��rɕe������y͎0н?	��I�SL���V/��-?����=x1؃a��L2"ڙ�G� �7�Yrf�?�X���6�b���d6�3_�_�
�m�2�����|�� ��;g{����<�+�S�B`����q{A��!F������}�z���6��Xy&{sD+`��'�����鱦ٿα����5�B�:�	5"��5�۵���>���?���RI嚔u��Y��ֱ�x}���E���u���mp6�9���$�]du����Q.f�5R�s8?����@!qJ�# ��_�_������`Y�
���	�� Ą���]��\Z2�nX�\��E���j�� 1�3�b���;�u���7�t#�������)>���V�1bQ�2����w��#��e�\�հ����,_�3Z*e���-�_9����}��������¨7���=2{Z��&�3��H"e�e2��nN]bl�V�嵉6�͞�P�!f-3�R��K2}4���,���޸#1nS�jK���]Hq�=�jfI~��e�#7^9ǈ��1�����=��K���W�I���(���������ϗM���#fL��(�h�%�FoL�X?m����(*|�Vj%:w�;x�3�G�c�$���xL[��=)b+�V��2yz�ȠW,��9*+�4� 9�ILԸW�� ������r�Ԃ�ٺ��3"�����㣶'�溆��󾺵e������{\��||-�y ��y��F�M�H"�|V9�Jy�bb�����#!���b��D��BZ� e��s���/�_N�m�����j����R�2� �j)�rβl4��~�yq���,W^O/H����<�T���F��=�/�H�:i: ��e����>�Q�{d4�z�=m=[fY���@ҟ[2b�4ت�vae�2�������=h�C�8�x���:cQ ^`����&���{�c3�5��'�ps��>���pv�걫��RVv��{w��ϟe?���|����R���)�k<�e�<@��-�&rDp���m��k]3v��Rʩ��ܑ���b
A����+�o�*c���������M�w[�����"�Rs3���k�������E*�ι��Le	cD
K�,��ʅ���4�j��fF�@Xs�C07�g��Jȍ5WWرB�f�����R���i9�1��������n������G�͑_�+��F�M>[��O0�z�c�s`��Ӫ�=]�	�M��E��Ԝ{^�]�N�sɢ�ݬ6���#��an�0�	��v9ɼ~v���Z�a�V�on�l<�d�K#��gHN%%E"��������b��F�0�Hi�k���'k�;粲�0�$1��Ē��������0���-�a�1�@�u-=o�x��&O& ��'�3�
1 i�`ZuJwt��>Gh�  � x�/�j�B�6ڙۑmƚ�|[���f�q�k�16��~��.�b%o��Z�߿s\�R��� �R���'S�6��� �>O�}i�G�V��;{���P���V��w]д���g5��s�O�!�?�{���3�$�gF0+�Ʋ~4y2Ej���l�:��#[3�G,b��]ۍ�Sk�<s�3���*�Ѿ-h����cQ{��Q�3 S����x��B�`P�9�){jbn�,%9*���+m��Gr���\� )�1�sT�� ��d%BY�~�@���X�n�*�~�ֵ���s��Q.�~Hv�J^2?>>p�0�������Bx���/ ���.A Җ���d�9恁2h��`��ׯ_�^��E_��E�s��d�ۭ���e�_`OT+���)8�q�d�������\����*6J2:�a��r/j�� �̂�������V�вl��?A$�hL-�G�)%3z�bj�3� ؛k�4٧'<�Q�%}��&4c��^_�+�ix��S7�no�=ڌ���%���	�O6m8Q]�`�F���F���=�������]���jI���\�kY�������U�4S�koޏ�?�;��Bտ��V�ZἯհ2q1��Q^_�<O=0k1���$}�{�6׌�ٳx��caL��� �|�<.oo���gy-8ɨ��M^�O���	�˂e�xߵ)�/K�o�5l�D_vst�R�s/�2���������ۊ��\ ���d�,��^#~mνD��fy�����3�1�(scp�h��VD�Z4���,X�����L�`�&���M��9��z��XN?ADٌ`�4�[G@l	��J1���>=ϒƴ 6�/��O���.);�}�bZ�9+N]kw/��g��g�d�����b����Ӈ��=��S�S,!3�/۱Ιyߕ����4J�V�V���v�RHBY�z,�#" +u��V���D���a˙QS@V��V�R���ϔњ4�G�{� Iy���­
2���z�2�X�V��H��yh�͌E��:��enoɆ�糩|Yr���r�ۏp��k�������e�{,��.2 �(+Y������?���o�d����c���C�9��t:"D��͊/���c�s���nQ�@f'͉"����uY�b?o�R�ǔp������3vn>��༯�v*�M샙b�p4+3�����fۓ�&8N����<�����9jV�=r>���9��� ���1�����aŎ�f���ו�V�uZ}�)"�>�3������75���h�xV2R\�+����?��Ox�H�g󞌾�;_����C�ޙ@�)�GcX�3瓼F����d�x�"\f��;���|ܞ���5�5꠳U�92��C�'ǏpNo���H�E}�8	�����zŏ?r����Ǐ\5(Q	������r)�.+��e�d�X��^/�����?��?!����7I!%��im% �Ucu��w�e��&R�����5dG^fMp�\����zE��l�-u�ey�����~�����7Ѷ6���n%��U��kDJm�@���2bƂ�li��dΑ���币D�[KF�,�a �T)�3�=����9����,�<�h�9v�� �Y���tu�����]�ԺRW�?V�u�(�����?�g��1�l"����:$ }�V�G�D�V�ժ��m� ����{Ky䟲�����{�k�GTϗ�xd�<KbJ����0�����/�%9x�)�Y���M�&ǆ����t�|�E	��ٓ%�ՠ0�:/'���0��%)pKn���Z��Q�������<.�1D��x���;bJX.����/5`�(����Y~����W����������y� �qx�	�C"2j������%TV4�������9�ǚ���۟�(��	P]�Ss�LY�n[>/)�'�!L�k6�#�.�R'���ܛ�\�w�\��lL*�� *�+7�Q~D�Y"'���d�4}n����쟖G�R������4K���n�(�)1�ٴ��ϭ�.F�6�ɍww]Cf�Ȩ�G�����$�f?x��Ϭ㏘��xm�R��ھk���̐�ຮSn	^�+��)M�SS7WŖK`��.ǫ�]'���e��fs��j�Y�*b� ���$)�I����Yl��t��X�`�m}��;:��x���<��8��&0$(����ʵX{����%�����q�����Q�ٜ�nx���T��J��[��n+.�>>np��q�Ք�:c����+a���]��e����z�ۏXo�[_"�7w<����G��,¿��������fز6@�aue���f����d���Ơ��<(��w5RkF��a@I�E:�I���@�CȂ�8A�7@s�q�O�`�w�__�s��l{��gΚ��R���I&�V��?�~�h&���'�|�4�w�H�`)A3��93m v�6 �Xl�X�~���HtόH6J�yƽ���;�n,����=�uO�,E�R�{`�b�Et��l����&W�+̞ޏz-�F��Q��=�܀}���Z���M�`��&�}Y�.���ᙹ\�/,K�4較�����ǯw��-�s�P��1_U��e����O���߿�gT^p6��q!E_M��3�J41l�ƹ�D�!ĝ���l�����vm��=��c�6%�_�����?���r$8�G��F�59���^�d�UDv�Y�yt�z-���̖*��^��>����?�Z�h�荻����ryȇT_㬒�}��5���g���C�����X�|��Z�@�h ��'�6j�{��N%Cj�ų�XhKa�YQ�k7L]�<�fjy���'�t0G֏�w�]'�yo�q�߉�O�L�;�7��g��<��w�6�>V^m.�1�.��Y��s9?w��9����t�\sњ�� ���R�7��r"�����O��?������L/˂�F$D$��}�&�lnZ�Nk$eWs�mJ����yN���I�Nﵻ�����I3g?-��{���+�{����&��z3��g����7C_��仚�Q���}��d�Rin� �#����n��b��cJg�#8C��{�S���ו ګ5��'U�m��,����j�ֺY!�6���!���yF;Z�B4��bfXL��Nf9;���<�ڗ��!QK&��{gvdE��n�<�|�vQyt�Ί��Ř�o��wb�F�����+����*��u�]��\��,
[����1�Ç�T^2]\�_�����/����o����.�K�w?����� 9²r�}BL%���w{G�(b�	���1�m+��*\,��9*��s[�˥ђ�^)3����v][��|�,��r�Y*�t�������G&�#�Rnx��ش�Z����X�?�{@�;����a$GZ����3�l�;��ˊ)G�m1��<�HX
�������F������Xi�Ff�ThY�ZhM�J��ta v
�t��V;��rm/���"�t���.?�5-�e_D.5�����N�����R���Ԋ6�K �LN�~�8Y�A�X ��IYy��D��6�����H)� ���jK��V� ���{ǌ�|Kv����J�=[���]CRL�E���msNI��]����4�o�֩�������� ���|��r����j$�Z�͝sXo9 � ���?g�o�d�2� _X�l�\��8�d���Z�h+��c�	�y,�ɝ��?�������~&��/����_���?�\/��/)i V��r���сj�$����pFD5���~��A{��$�¨4��O�L��y��^���(U�%QM��켯y�k�p}�<b�zD�g`9���{����<k&�%����Xe�!��+�;י��wR���[$�G���*,´�w!��2���gb�cUT���L�G���ڕf�g���������`��d޳Y�mkc��`)i��z���#�^0�g��Tj�5[?�~����B+��Q�}5~De��@���^��-9��r�dй\�~y��ZJM���Q�q�De�H1�.��򲲒�˟����/��O���]�\���������$�A� �yX�Grь䲄k�Q�O�~_|?�K;�G�N�Z#�/dn�>��^�vmV�ϴh��f4���e�׋��5���;�}�"{�|&p�b�!�;-�\�"�Ky.3@ҿ�@�^���,�d%eBo*���1���0��1E��;̮��h`�{}�0�gB�k6�M�!�а�ܖ|���Rcu�&�m,��vsm�o�ߍ�B��:�˽�V;#F��kʑ��w�=�گ���G��㌙u��X	�1��W��zV	����[ۭT@{����{�V�G�x�=kv����u�����{x��㳿%W��.�lH@�F��N�Eb���do=+/� 0�Ln��D���'E; Qf
 8�Q�TJE�`a�㉟�7y-��^�n�Զ��t�Vs�Y � �\��M�x�~�ϱ�&�waScG7�!&��H$7�T6z>Vo:A�u);��ʽF��lD�X�d�3ɻ� ��N�<�$��?$�^���so2_��c���S[i���Lh# ����
J��S
����X��P�a����_V�P�~Ը���
9����K:+�>���36V6gۻk��<��ok<�@JO��������vu࿥IZ+��|d�f�u���X�#�5���y��k��?u}�L�:Uљ�r�����s��Hsk<��N1��b���$��Rfs��T�'����V��~�������%/����~��O���7�o��֜3!*8'8��$'F@D@J�>>WNo�Z�)��$����=�eQfJo�w����n��n��taEY�`�����P��~��/�ۋ������:�b/-�9Z�|;��n���'Ǵ���Y�ŪI��y�����To#��J���#��\lņe��a��ðF�e$��Д�ۼ�ͣwrSi@� �N�g@^�tН�;��J��)�,���s>\�9F �>��q#�����q���u�k|j�߹sn(l�N���_��G��g˲4����6k�ʗ�c~��ho>��.y<g������X�{&" �|��;������yҏ���뱢��Xk���@���,����
Ė��s�����<���O*��s�������칑�r�Snf͞���杄mo��<IҬ�Z�I>�r?���~{{���D��縑����,xs�Hr&��7�zA*`:����wYDN��Rf/S�sk��"+	9��y2�x����Op��\��;�w�4y�^��)�Ht���B�rT/kN��CpnY��=fv��rt�/����k�gE�j�NN�#1�Ԟϥa&�� ���W��ɶ��oh��mf�"7�8�Io���={�Q�|N1�܏���Nc�({m��p`l�R��d��n�����)�z�ܴ��gL�H�}Q��
і��m�`=��;`�m�fhw��5�c�ÞY}��ܪ�c�RX��ơ4�k�x���g�4?�v
���Du�#S�Ֆ��R�4곢G���#��*i��>��� {�D�ɼM���}�
l�S��*�r���M�'����7�l�����%�.�,Yr����"��o��b'���^�����"!z���9���"B��r���x���|��d�����w���c����?�3~��_��C���Q�`n0Z�F�Ƞ��T�f5?CX��Z�l��g�X>� ��4�X,@?p���,���3:/���T��Rd>���sY����#�]:�����KZ���&W�I�ŘIQuFt�w*���l2k�g7;�5/7S�L����y��\%`�ʃ�)�}睊��a`��&a���}ٙ���3�yĄ�stݔ6��4Y�I?c}�l"��tf��R׍҆����3�Us�Z�k��g����/r>�cJd��͊&�	��Dq��Q�Z6s�$��<�1%�k 
�Y�ۢhr��r�>C�����.8kz#@+��1�>nS��+�u �9,~�Y�?�wx���D����.��nq+�%�T��eY�b�����1O��똯+BX��k@����G����mF��ͫi]�*G�d���̭=fB����6}��pR\n�w���ϊn����X�f��'�gN]W����N��@���H�1��!�Fq�����ͺX}�@Z�Q����1����X۵U��+�H+݌9fc[�����tU���$鲽�(򞉶(g�}u3豈�y_=���r�b��.�����%��+�{50�s/G��-Hma"W��H׃B���2��\��h��ʏ����v�����z��Bo�,�Aa�R�d��jz��}��?+}# )�֬����Y%�����!���@����Z71����LF
���>&(d�E�+9gF�g���,�6��;����-R{�=�)u���hѓ�4���|�� 7]��'��V;=�癢�B�	P돦�wĴ������.�
i0�L3���b0R�_'xD�h��gG�|�#%��Ҿ�ҕ��l��J���:+�f��V�I1~���I�K��� �<�ͥE������� ���;�Hj���F2h�f�յ���o����h�TZ��gg�`Ǧ�1"��X��T�R�+eB+A���5-�����Z�҅��mU�����,qOyef3��~:�<߶�'~N�"�u�ò,5;?��`�5���#����^/X߷w��7Đ����*��11���\I�XXbGp!W�!�"@�c�����k��}����l3��,�@)ôF8A�!&B��|A��ɒ���ߚ�_�.�<�y$�� 2�N��s�~T��9�>�����|-�l�drF�<�	�0M�L��N`�;]��Y�|-zs���� ��9���s<����ǈg"M����;����Qd�4+)V`Q`����)M��A@�w���S��_�������T�j��������.������2 o�\����� It���J���2�	Y����Ţ��5���R�ĞF�,�`u9PjY<�GNc��j@XW����+�L&(�-�8�JI��?�3�Ͽ��,��S��k��{d��ۈ�i���Z�z,$k�5wft�J?Z��ڬ� }��iKf�_�L.�e�Z�k�s>S,��g���}a "-٧+6��z�x�H/0H[04�w)�������?��f��+�MW����}s���֊�̻��h<�-E����V����=��G��9u�(,1��]�Y��{�UF�L���`�w��$�&�'���7��Pb��҄v����]煍���M>4�O���=�J.̜�ݗ�)��*�0��Љ���,�d,m����/aoƮ��/*x��k�w���x�� �)H��	���?@f~�Y�oW�O������ל��-��~F.���x����;)r�R4�}F.*��Y|�!e@)I���3��V�h���Gb=�ަ{Vd��y�r���$8�Uph~����+�$k�S��J_���9����h��Nd?�>�v�s��V��X^f�8�zOs�A�]d��{��덵i;,�k��-��^�����O���GD�X<�si��`N�!��e�f
�\Z��n5�-��"Z,E>�PS��d���w� [�S=�_�'P�X�Z��2YT��bĺ�0VV��
Km ���q��N��נB�#aӹGv�sDa�~��ɸcN����� �UH��Jb�8;�&�9�ִ"�eB	�I���H=�!&·%��˒��yr5�(�7J������ҲCJ�������x��vr_�Ϧ�@
���7sI��S��1��s��;�\�T�z�<Ϻf�-�Ge��{ Ќ���=}�a���u�u����vy��	�~ͳ��/�SR��է�}��4�8�-�Lc�Q�e��aN�u5P�{�ز�Me_z�jK�~'�{���IQ>�#`�?S�Se����C\W�!���4��#˅���P�\m����(a��Ǟ̬�M(�X�w��t{�ZӸ�/�6{�@��v�кm�\��uFk�lj���1����Lc��y�T�./��d�5��s���F����W����	n�RL���6�GI���׈A��RbU�����c"���-�e DcƔ�{6�n ��D�T�y��h^LF;��yo�g	���������D��f����@�g�2���?G�1y��PF̘�
��(j�T�߱�V��>���̀9��i0t/�.����HHl�^:�˫�d��j��݇~���]����n�Υ�i�Qc��Yvڔ�g��3ʞ��3��{��{D>#��BIf�Vz��=�z6z�.�GJ�U�W�u�d0�x�>��d��
v����Qn�G�cV<`w�G�;�%2��䀟5������Ļ����*�5���R�@����?a��b�!3���w��\*�#q�v+�,�����W= ��|��MV��&W}bJp ���J�ir�֦򏡁�3�=Y�d x;x�ً���6�������N�}���eXY�ZM��G�JDތ�~E�;��ӿ���Bτz6'��<�~��d��9�u���<b�>�IH��;���+�vr{� �m���c������
Hr��j�S��g��G~�R��2š�?�s�U�:�`�T�j�"�<��jf��\�f���ne�3�uLf�%�%a3S��DX.�5R� "�H�A�� #�FD$j�fS�N��ڶ��"�.��hK_�~���zg"lҺߚ���iy���Lq�����=aC�����]I<"�J�>�i�0"�<�.`Z���Z����ygX6ݦu�#L|L�7q�:��l�,���Z�jXϱ�S�������
M����^r��ycϜ���sή�=�R�?�<�=v���<{�xGp`�2F�jnO�{ޟ��G�t�ҕR�n ���sp�֤~��- �y��R��/���3ƈ[���ٺ�M���"���\�b�pI��0����F9���vCX#��˖��GBk�p�4;=�����jN�$���]y�]wQ���o���|c�5ܙ�~#��;|O�����Q
��F��7̓/����Y�~wg ��yt�ӛ��%E�)���}�S��g�/˧m��HH�iFF�ov�.�E�5���^�2{i6��)�fSI%�y)]+�(��Ɔb�v���VO���5���w�ܨ=�:�B���+���	����T�X�c[K�>���_>�M���T>�D��n��.���VS,��4f���I���D�a�u!<�_pY.�u���!d�Q^_R���nXW�,������י˓P���' (3G&�A`�; ��H@$d��rlmE�M�:� ��L��{��z}�iM4��cc��?L��޼V�������jj�yf�g�g�{�d2��'�Iқte'�8���$�"M�s�`����vՌ�xYg��U䠹�� {�����i{ET�x����6�J@�U$Sv������˞�@�g��,�	��Ƴ����ו��Yb���+p��d$��4�]�|��ݺ�-������O��<дޑ^�?�ۈ1��><�:D�p�|u�C��.˂K!�����늏��8LfP"�� p�$ᫀ�Wk��`�0� ?�,Տ1��z��$��]+-�=��{׀G� Ejt ���ED,���g%��*�ґ�w���(VE���O~>\�(v��^ �).Ks����� ��~�@�g���f��3�������w�g�_�F�^W2�Z��9__�^�5���]��(j���#)�d�׹89v ط�q�)ڏR;)m)���g��k�G����Ǔ؏H�E����˟K
#�9�������������q�5?K^2���@�⢙��ʸ��C2e3���њ�U�B�V,�q�֏�ݷ��3m�8N{���-�4U��*����zVZ%�W��E�^'m;���c��,5}��`��f���li��a���Ѳ�RB
m�g$�>s~�Iп�:��s䱀(�-��Zs�]m�)�8�o�Y�}�߳�C�M�c��H��͒��]�֚{��%'(��R�:9z"׀H��ycG>����κ����(׮t�����b\�}@��{�19Ҭ��#M./5愛�T�)!�X��;���6�9��9Py���W�k}2�4��f"kS����	K"�����p	) "�3�#��^�0wUv�x��u����ّ�W����G�Z�>u�o%=�@���EJ�"@z�H/�%HhtU����_�$5 �n47^<�##��m�Z��N���Ə��>@ ��֔�Ww��Tc�G���$�AP3:5�W1�@ay";��R4I�+}[�Yv�{G��$I�N�(�RL-�r.-3��&h��pY�K���՞����?*ԖU�q&�R�p͔V݃r��<�#р����dzઙڨ�7r�f�	�dc <@ÿ�r�ڸ`Y(�_�>� ��i��}$�c�ܨ�w8��<�gsVZ��� ��d)#�(��d_�Y1������Y�ht�}b.%�䁠�l��e�&%�o��S*�$`�l(���Y��qM���yc��e_
%����!����Z�eIk亮%3��`��3���~���{��bA��o���&7@���?>>�?��4�6�����{_��w�����=�ł�ŗ���4��w�s�p��f�G���3EP����ib�ބR��rg��A���sL�1���7����:��l�Z�cy_��u^����g�d�E�|~��,Boa�Xk+�0�|.�,�ϊLέ'^��Ԓ�V�=��Ro��R{R��� q���ţ��J<'��w�0:�<<&�v_:�ߑ�|�g�̃&5P�mp��ָ"��k�Y[�+��fǫ���Iѽ�\�/N������M �i����.YO��A؍9���l<��6#}�k�ɾ����}I�S�5D����d����@f4���f�[L ��D> "�,7���&��t���ś�)ڮߖ�ǫp�1���c�����Y��f����ru��zy=���� �d��F���*y40DV�y�iY2��f��@B9��e+�I�
��?��zFv�<��굞�o����$Ư�u�h�bk!�,?��ӓ|��Y��2���<c�Z�<%P����J�y���X�WM~����Q�%}�R2r�*Ĺ\A�:��u'��ފ��uML���V<#o�튘����9�<FD�B!d��&*�Y��ڏ1~���4�p���?�&�)9�xD!��v�j�&<OMhzke����Ѥ�5aj�j��3��-`�̳�U��Չ1ZL��\܊��6�2�j�Z�8�c��^�����\R2gcv92������ə����3sl�3:���鳑eC�Ƴ�dD��mc[ֻ������<,u���3�ƒ�<��g�&�r�\/d�s)�R��t�O��+q�����K^#�L�y+�r��W�>#��c �a �М�>�#8�l�ǚ�fmN��^B̅`Cb��������E`4�����^E�T�D��>6��gLJ���-B8ɱ��V&Ok�Y��{�s�.�H�G���^�D���g��;���Y��gD�[-�j��\�9���lE��>o�ܚ�ڳ� �ֹ{��'�t�����U��:+`k����u~O�mF��5H;�eV	ׇ1�]�7P����n��*C��+|��o��ybT��DW�_�]_���Ri��*�m~��͟}�j��S	�u�U����C��=N��v��<��6�k�kr��a�+��z]R��\�:�n�P*:�����n�~$���!$���o�ع��q[����Db�@�*Q"L�tFؑ�Ix�kw�ƚ!W��Ɓ�:�
2��'���_�|�v�H?.?���41�������[&n^|Df�Ŗr��&D���*�ѩ�*S�tկ`����ѱ!�Z^�dJ_��������t?�͒X>W�!�?��g�V�v��� ~��|�]�
0MHjm
ֹ�n�z�b��;8ld�.=�*� ��|"�m	7���/1�d�֫Pc�ºmz���K���<	@S4���zI��A&{kC���'>��ۯ_p�vƛw��|2C�C��d8!$��
 l���@�[~�hA�w�إbj�h��l�GI����0+����Z��G��1��*b�qlGLנ���c^�}��Uo8r-����|�D�S?�=@�|X��|�M�hJ�5�g�էc�FB�c볙����h&��.�_�ko�.�w\� I���m��k���w�h��J��*�43��=�w��\G��y@�cR֯er�5�dsț�l����[X;���*_��� ������cLel-�RV�q���1�:CU���ϊK��&o��BΧ�Y�����v�R�y}L�;�p=��[�yL�Tb���{z�m��"�'4�C����ᓟ��K�ڲ+ݷ/����9*R9K_��,Y�aڥr ���g�h��Ͽ�j �L��ߓb�X�G��>�^w����z83V5YaBq�ST��:���gJ�_�����K�5�l}>;ofL�\$h�~�3��4�z�]�"'���Dys��ns{�����P<��c���\��Ot�GdY�]0%[������e��sP���0]�y�\Ki�R�BD\��>x�O�	�1�$�H n.��	x���g@@��Z\��{f",�g>�\ұk*�D��\ş�l;������s��>�ٰ W�ZE�O�SJ��--�I���^�pu�0SWs�򜹺�܌R�'�Kg!��-A_��4f�lZ���%��K��ұ= պ��k�7)�>g�0�#�92����gg�]����Ym3�f��2����'�'��L��'ȿ��F�s��m���S��.`}3�f�DJ*��'�2������l��G��#�s��+��8��^J�Ѿjs��>:&�r�R�=qj܇��S�%i�cMc��a-���O�0��a���S;�~�*�||�v���:����{�1�V�`a��JPZC�(��"c�Yaq��:�8��Y�M�@Nc��K��o>�E��Xb��>�\2�� &��c̟G�~MlT�XMz�\�:��E��\*�d��D�G��P3x��ASO*U>��6� ���'���G�B�i����w�|�Ll��F��d�5��RU����Nw$;��O�� &7���$��a��L��<���*)���F�Ů�l�2˦N???�c��?�`�f�*���yu��WKk~���oY[f��b{א���m�]�9G�vk�Zv��D��Z�s�I)�$,1Q�SNPP[��v0O�%of{>�gH�y��	 �k��\�_�b�9[Kn %��:8k�ú��;o�������W�ܿ��1�<��)�q[�k�y��'�2��������▔���s|q1��-.KN'�}Π�֋/7]��XA*��R�JR9��������qu��h�׋��h��xvGΕ��h�߹�� �錌��w�ƴ����؛� �Ǔ�̼���#��ڞ9����5e;|#;�<�	����$[�mR��	Q�3�d�l���l۳m�/�m��Q��z �h��1n�ҍaY�u�ր�]Q�K!/,J�鳩x�&Ac5�_G@&O�M�!��k�}i��d�l/DB%��}<ݒ �u音X.�5�~@&�r�@������u�)�.�!�0�����8����� ��Ah��%�k�F�J	�24м�&� ��l��-��D�&���yф
�9�2 �:=e���2�)�n{|�Od:��ot/��Mܴb�ϴ|E�����h��@$}���{,����'��j�syd�:Z��-2�9���H��VN�V��V�ɧ���K�tv��Wn���H��<������v$������m�f�š���EoK?���h��\�fE�����\-X�=�PGuo�j�I?�1L�E}���{_y���m�d{/�ӷz��g_�z�[p1�¾߷5>y�=��:(�N�'O <Y�RG2uR՟<vW�5�������Od�#�t:1"�d�.��,�	:y`�dJ�1�bӭѫ[���T��\�wf�����Oc�,�RVr&�.Ĕs��-�é��h�S��u��$�$�) ���8	�4β(#d��E�X�Q�^x�FJ�RBf�J׎� )���ψu����6$��#ُXn�q$�{l��%7��g�k�'1]r�Ŷ?"?���V�x.G�<N��P��z�<�e�$ٯ��`��{�˟T�O�g��g�Y&~vI���?�u���um:����q�lC��(�kF�,�;�'�ӵ�8�`���*��Bf$y�I`o+���Jk��/n��m�ucM�IZ��=�l��Y�J�A��?���69,ˊe�`Y���3G��-(��,�#l�/
|��|'>bqnqp�������5fw�?Ā<B�F���m ��%@#L �gI��&������k�X�G�[��|4���5��e��^v�1�6��`�$H��a�)A(#��Ǭ��!-s�N�v@���s��Z8䎯��hʷ(�X��DY$F�� �#f�wJy6�oRfG�m���=�����?#�l�TBG����|%:��1��2���ǽA��g�h>"3�G�����ƣ2˨j�G�,��<	 %pܻ���3��|�y*��Sv��$�d�jg�Lx���|�0���<ѻ�ybx�؈1n��,ӹ�~93�ӱ֘3�@���^U�0!�%����纼�'3W�At9�E�gsy1��	=3�!&j� d���Kf��H��Tu 1����w�	MF
j1�(I��9:�8g�v�g�eʹ' �g�v��b�j�7�#��G�}���#� �#�ct���gۑ�/��z�%�� L���Ôr����fE��ƀc�\.�n�
z aY��(���ؽRzL��}��(�C�m�W���B�')���K�F�T�.�e�%݈����3�.P=���W�����ul�# �M��ͭ/�� ���LJآ˓���sι��>��<�\��:��,�1"��8�
����o2ߖ�3M^$syh�����T�����3���|�0<�����1�� �9�>�۬P�K�!�T���{��^���8���c�G
H�L������9h��-�
�TƲ��'�{�W�_a��u����Z�y(�#�c�?��� ���jJ��-*���ѿ������<��1���}�X ���L*��Ti��f�����$3,lo,������l�.�S�;��� �M���%��?�8���wA�����ҭRd�M�C���|ą&Ϭ��p�G,���������}s��)�w]}�_�T2��У�7�k���V���Z � �e����R�
2ӧr��?'%�.��O������|b�����ֲ�@e�Y(�sH�4(Ч�OO��dF6@̓"��)�<�n�eq	U+��{�"�C�u�������.���7� nͦI�,�s{r����ұ{�Uo����w��R�v�nE�s�ghu���,���ia��(�Τat��CM�@��*`���ԞO1Gv�S�Lf�x�4{Y#vJ2�_�szm��o�X��{�������g��z�,��������$(zV��J\KJh�������#���{��C�R�*���q���҄��<��u�ԕ{`"�����՚��il�9�����i��&1�������d�zr��'���q-���~�}_/x�w��<�daA<3u�Nr9F�SL��{���izjh�y��Ѵ�:gr�������ԧ�fg�������~&(AH!�d�vHh Ƹ���~�T��-,�+�(�s���LX�q>Fa�n������o�����ԋ�m ���"J� ��j�,g����nƸ q�2ƈ�PE��	d73q}������̟��i�GQP��F�
�a?[}E�jׯ����-_�g{	�R.��ߺ]i^�"�����~��&m!��3��+.#s�3�zv��}ڝ�E5��5�#��̇��m�\j�������ǯ��ր�6���W�/y��F뫤5����&�3����,�lS�];F^k�	/�ǘS�lV��.mXIYd�@�2>��N��H��m���Dݔ�d��.����@���X4�&ͻ_q��\�w�`P�_&�a�\�����_�q]c�7 �w �{ ���M}����4&��)�'������$p�Kz <BL��}�� h�r�r��l��3�K��:W��;�mjm*�kxF�).!��zv����r�Ak�WȜ�ܥ8���x����{�{��<��m�q*H����!�"�/��8�=�� �/�2��}��!nf��g�O�l�]ü�Ҭ|oR����3D3�j,e��Ez}x他H�*<>@cwgH.2��Yn�J�al RZ(���g���L����gs�$Sq�?"�9;��w�u�>���6b�e �2�ܽ�����
�,[���G���5`�� �oO��	�F��쇙Y���h3�'`����3����	�/MJ��#(��HQ�-s�^��I06;֩ua�>�dRdJ�ٝ��?��<l��fGKۢ�����\elv���Ao˼M��Yו9y�
���i}�= +gI�I9�e�e�)=�d��z�4_����pT�b���k,�Y՗Zօ���&AX���y���V��+�z�J�fu5�G~��vW�*�XEu�6�x�I��#����z<`��k�3<#s��X�I�6Y�%�,εa�䂌�Ɍ~I�|�� ؈�F���7O�Љ�F.��%�z�>d��3f��"ʷ$�i�l�C@O�j��&Pi �sp˂�-X�1�S^Np�=��|Ȟ1�uT�G��k���2�����
$Z
�=#s �5�K2���j�~z`��<�NʌI����fLX�h��4�u�����r�|$a��~�6TaΕD峌j��(��g#�5`����1�0̇�ۧ���Y��M_��-A�I���-L�am�!�T�v:�ƫ4ӎ��M�yP-��?�o���~�\s��dr�cJ�~/�����^?RC
v���ocfju�b �楕털�Z�J={��`~\>R��J�RT8������ӫ�&����O��ԯώ����t�R���0�|�˂k�FxY.	_�c���o~�.�_���ZA���'�XI���JQ���D��<�0�������# ��T��&%�@6-��=+i����~?��z��⬍mW�����ra��#ƀ T�"�J���+�~Da%�pS������+��cܙN9�m2�<[Cܒ�SD�����Z]� �-������lT.�x���c����l��F�u��~���P�yk��IϢ#?��x���?s΂�Af����)��U9��)^f��<��]��'�v�8*�������}���v��H��`k�,�<���LA�_rs�<�&�Fl�7,	p�hr2���E�H���r
i'�� �W&!D8�*p������zk�ys�32���a)83X � ^g'�>[I��g�� ��k���>*����A�Ǩ͔u��砭W?�]�����2��y����-٦�0?O:n�F="��Vu滞H��1�Z�ɍ!�[~fXU~\�^T�҃��ڍ���ԇT}-�X�L:C���@���~N��;��0��Npx�	��a���!��L95�u@��P�7G�m��������%��V����%�\1�o��i�5"�|ҕC�Rr���X 	���Fu�L�K�E����<��� ]�ZW�� Tʳ$q�|A�[������\-�jg]�����y���e�y����Qy%���ӡ:ڬ��2|���g-Vb���[mH6 Ư�f���K�.h6�_���\6|��u:�����bI�1����gsg-S�-�+r�BI#t���H��P�kJ)D�Y�X�e�ā�k��cf�%��+� Z�I���?��g�M&;o�\�X�< �d*O~� Ȑ��)��G_@f1���C�sor	&=okഈ���1��y��0L��Y8M L �B�h�N,hi꾵$���ˬ�����-�~��n���o۱��A=��w��� ����8�V�:/$��,[~Y=%��L���he��Z&�V�~���f�b�}��w�+O�$ �Q���#�Y��x&�JG�|(�u�'40��(X,��A�G��k5�I����=��^��,�Nc�y���K�M�X}s-��Y�ƣ�cL��u]+�9������ȶZs��_��=�f�j�ԉ���Θº�s4�DQx�f��)�ד�ү+��kmUf�
ء�k��=%��6�K�˻�c���{�aw��\��2���~��ki��i�����xʫ��6�`{�8C���e��h3Wi����`,�����cI#h���w�LD�l/��,��l.�u���"=Db2A�M��&(����2y�C>?? �-pn�E�I�9b-	<��ìoN/y0)֔��83������}w�(��͟�d2�~Lf�ip	��C+�6]g���;��&j��F%��m��>��P��
��1͟�}ڀ�����j��b`���*����X7��3m�ɷ�ld�ԧnp�������-��:�+�I)��]O:c��89�,Q� �WpJ뮇s����ڢҐ峝�c̨��@�r��5!�d��r.�aY��vY���|��/�Q��&'tft�f"��E�w��@7��Dh�\��٧]O.{(w��$����l��ؘmrP��#&�#��I(�h2��B�Ǹ�y���ʮ�O�_=6h�b���JGD�4�������[��ʋ*�P�F
��c\�k̊f)�m�0�R��<|�9�WD��ٱ�*wɯ1��c�?�uz:{�ld]f��6�a���'r�K˂<���蹚�Ck�u\�|̤�Ef8��X���&�Eb���
�,��X��'��O}�܇R���qV�o9.F:50l���������~/ ��,�{q4��p�j�R�۽�\�Ε�T�ܘ�KL��\�8���=����|���\�#��$�u��oM��:�1�L5�)��`'y�)@h?<�MZ:�H��#����d@cʑɝ�S���]�y�L ȕ���L�e"Z��, k�᏶ג����L�g3�#�q湏�|�jsa��I$?s�G�'���v�z������`�]��$ۦ�=�{�����	�!ƒ���o`?i]"�v�u��(-W1�BdȜ��c9@$G^.9��Ur�x�k:�S�GT�d�@��I�O���=�~��S�s�s�s_�x+$R̉m͈���ls��}�ǹ���p�+n+}'y#��=�d�?)&�az��'3��b&P�o�F���1�ǈ@��a�(���şbd��n��cq�^S�C(��"R�����nu�s�D��ץ�������Y��?%l��f�q-�@(~,�;W���Rf��Yn�1;�{f��g����F�#F@s�0�����wY9��8�,g9����d�۩��V��v�0��h�h�{~��w�򓌱J.N�J4[�ִ����?���]Ue��{9�=��D�� ƖV����V�EcԯGd�N>�����&` U��*���?G`j�.h����΋֥�矟��\�U|��L�<����l(�I�9�6ܲY�.`2�|����611�?~���z��w�������;~��_q��p��Jۗ˲+�<��b� ��h7Kղ,�5%G�}]�����di����1�!�P��(�|��_Y=s��(�Ɍd+�힭M�l��И��f�GSq�b���!�{��f���G΂M���YLjs���s���}�T�&'�G��(�5-�!٣����y��3����d��_����� g�ؑ��d��/O�4 a`4���]���"눓��`�@����^��@"��;�yyP�\��W�Dk�=x�"l��5�I<k�o��^h-��5yYBخs��oW�[/5�Ƹo���a�����W�L}y��<���X�|�%�<l�2{�4�'4c�"K5I}O�ky��.��������ܺ��@V�9[Zi�f�C<"nG��32�r̂�3|������G��RɌ"�k��Y!6S�^��&���G�����r�'s���3 L��kw�����eZ�/�p�y����Y�Vn��F��+��l~�c0�=�tsG�S�=F2�?����Q'�Ց�Y�rH�zt���o� �\�av�Kˡ��6X�˓b4��b��&O�u^|1CʍY�u>h�ؘ�Y�����SU��N����
�+�~^���u�d0e-�R椔��$��"���4D�d��=��i]���x�i���3�96@w+�e5v
����̵8˹�73X��Z��=�)��Lţ�X~���/���-dY�2tT8P�r�=k��8S��|�Zl�|>����g��t�R��Ȝ+-a��!n���k�K��^һRXԃ�k]7lB��i���J���XcsD����Z�2��Y�D����lN��̲�X@���ؙ/f��Sq��s����d �ɩ����`#�aR-O�C��h�1Z�N�1�>�:�<ƈ��O�������?���Ue��^��.�5���t��� ��r��s�n�`�G�T�~Q�h���Y�6�u<�]����,�s��C��l��gڬ�3�W�Ц��n�Z��z4�|0Ÿ�m���+���}� �|7�}J� �Y�Z���=�b}�/��6KZ�΍��G�e�h}���Y@ˏ�1?ʖ��4��,B���H����]�N��s�, ����+���kU��E�,�i��m��Y8��8n�l��ٸ�%��1��>S� �X���n+�w��.�k�<
}~~w���`�>`��" E��˵<sc��O;`�8\��|�\p�{���O���_��	 1�1�I}�i�|���T'_��rB�	T��(r.6�M^�FSj��x�A�1���#�3--!)Zo�����WW8�1�?���ئ�qx���Qi2�/`�%��K8?ۗjv�4�����e�6�Z���2zo<5�+�]�?�ϵ�8'p�A�3�>��DK�C�}a��F�W�%@/���h��z^-�������w-�|ؽ/L�����2���JI�r�MV
c,@s֦��>?�R������1dw�1�x�Sv��-��ߘL @N]��;V�Z~�9'W�LTz�P�`>�_��Q~/�O����恵�]C���W��H}�x��m�8�].�?��G�|�simF�2k���3�۬M�J��29�X�V��+KMr�X�:R�s��D��)��ӳ�������>����:�J�#G)�4�����,�q$�e}�F��M�k"g3c�p."���1��6峤�b]S��RZ2w�8��A�������@�5���-��~<u�g�������y��.�����=�	��2��=J�zm��+�����N�
����$�����,��ڙ�.^��\�i��Ib�jt���=r�kπ�l:s��o���Dj&_�t�$��Ϫ=�;�ɢG��3Lgl?*`R����85��%��u�1��
��y�y�Ej����ذΕ��=ؘ�ݜ����|�H&|V?�σ�?�8���q-�}�����9$�G�S9ɐ�j��p�|�4�I��df�C�Q�>']��>���k�8*�҈���1{A@����4x��S����R��zE����+[��E���>ɖ���g��?"G@����`E�&��
̲+#E��Y���w��Ҕ�L����Ѯ��k����)�Q��A��Sʭy�U�*#�\�  k�6���ZĆ��2��,�:�r�-�dmV��}s�5�\��T좔ݳ;�v����y��9�Ffʣқ�{S��ye��c(��i~�#�Gs���Y� i��g(#�վ1�L5ϵ9qd���W������1����ʐ���u��D�[ �:�~Y.�R��C�u�- @��eqX�1n5��\�\	f��+.c#>o��!`���[ޗ��'S���d2_����k���@��{`��Ofir�SSM�9����g�Li=��u(�Iݛ�9��8�ިT��b����!�����I�x*[q�*��l�U ��B����2�7��j7%�HI�4#��`��&ږ�������s��K��K�۞ٟ��F�l�^��5�>�/Fdû��G	���f۠s�|͙�,	��_��Z��e ���[�}c2��|��,@3/T'���x����1���*i�WO~B�|WԮe~Q�6[r�y�����=��h�*��J���qƸEl�k����,S�����>�@�W-�;�j§��7D�]L�� Q�r l*���Aa�ZL�����7�����k�e1_-=v�U���������3%��4��M�x���m�1�G��;7&|ݞ���X�
�ሥk��#E��Ua8�l�>=���<W2�¹�:�՞��j�ĸEo����*��1��C,���)�'b��r�����H�;F��ٕ޻�w�ڱ:���r��+��B"�}e~��Y	Ky�J����+���i��5J�������j�y��1Ƈk���V�n�(4�g�Q��wb����.ϼo9�~���y��v}�\�[j�����>e�e/{+Y�'�̷��_�yU *x���2�]�50qn�j�
�
��6>ƒ�ׇ2��r���`���O\/?���K�m ��o��?q�b�߱���k6��Tr�,�1��1AM���6#P�� ��$E���9�R=s��I�z�֘�%R�Yʙ�`����P��ߌ�^�|V��>�R���\����~1�����9�{͚��{��<rMfQa+���L�0lm6����E�]8)�^��#rT��^g�Pq�0 �]��F������x�����A��ٶ帠ϸϦ��Y0������}�f�������ݴ�l{�?|>I�rO��'��cSی�x%��%'Ɣ�������ƚ��M�M=�7�w4c�=�2�o���2� ݣ�a-�f���3�qҸ/y��}��k�U~_��s�䱛��M�!�䀳.��g��5�養D0�pa��3	��z3B�|�	�d��?q��p��F	df,ҿ���w鰼�4Q������ �����!�wz"t�d��Ѩ�#����`P6�h���|u�KR�j��<?�?���:�O�甅�*���"�gM�73�� �W>Sٗ�Y���bL��~�g�s@��>[����l��dlZ�X�9�odE�=ପ���.4l��{�Vk�KZw���J�'�rYr*�t��v+�Y쭫ɔ�}���~-�d�,�����ؘ
��`��W�[�J��E?.c�ډ�SnM�$ɟ�d�M�vzȻ�Kޝ�J9��8b��Qi��?2�ОMI��
��z����Q��L{��R��ʤ &�Y�����g�+p�<��>�G�?u����f�?�/�z�#����8�{F/H�6Z�����=I���wHY}�˙���=T+��k�  �.�rg�R�'��|�6��$�i�IVX���uָ֩�쾵)H�-KJi�E���6���W���;!�d�f�ʶ�LJ����l��H���r�eI�H!ŏ��`dr	��v��u߿>��;E��|40h�����z�史˚ɧ,��6Ki�g����p�SxpS�6?�i��7S�G�Y=P1k<�G�V�ܞR����%ޗG�ˌ��YC�9y-���-���U��쌊g�k�[g�3Ōl$T_��޴�t��2_'���֚T�fݛ��P��?�&u�瓉 �誤x�,�A\�i����"3�t]�m�a`��b��ߟ.\/\�\�םI4�������/3ƀI9-����v����ܲ]��Z���F�7+OJO��$�r8e;q� $�"Dl���[����H4-~/�ؖ9�[�����f���;�1�k������գ筙��ʹ<ۿ���|V�Nsm��)���5�����H�����`V���˟\������҃�{+ޕ�Zc��Ɍ���>��Q�3���ϸ���T����X�K�P��ݲ�Zk3Ԓ�?����� �d^_\n���)C�U����P̖�����Y���=ZV�E�>��C�S�?
�L83����/�1����$���BIk�,Ka2ݲ��nY���ʖrۨp,0��5JK��v�G@�E�@S�G�8G��Q9��h��ߴ#��[�^#�mc�A�,�y5h�J9���5}�z�F�ڝi����>�����1h����̿��
t�+ףb̖�X�>Д	ٟ�.�:�i���E��GR@/�o���+'��㎈��nyȌ)�H@67Ƕi<�=l�ٴ  RXB{�L%M��'�{_�����+=�k��G}2�^���2�G�45`c��.�DS��j.Gnk��m����}z�.������2�a�Y�#K�{�p���J��g��?��ќyvN�}��^���xd.$AxK���@���ԀJ;~�3RX��3�\>ǔn�D�/[?�O`���!� �~e>:��E����@i~� ZJ�j���0�p	!b�خ����3�n��
��=7��ZdR��hNؚh����3��E��X�2�U�=�Q�(C���yE��K�őכ� :�[�3�%3��C�>�7�UՊF"� �"��Ci��D��g�qO1{�d�B9�yj���~V�s.}<�gY܎���>y<��1��v�����N�՚�1D��b*��M/��G�����G�%�5�?):6&�R6;F3OS��w@�Ir�vX��v����g��e�/�ƈ��O\��M��{�X��=�����c��%�g\C
����a���#��
�(���wfoN6�ᩝc��\W)(�t+�Ҿ�L�dm��-W��х��4޾&-����������wN�����g@͌�6Z���9��T7�G�]$�Xj�S���G���3&eR�ۃ�Z��s���g~tj3��Ӟ�]ymy��d����޽�Ha�}|�\6��^��f���L�1Ċ���U�p���G�
h�[���lKV����v���m ��wkY8r�����oV�����& ��O �0�$�ʐS^�u��3n�3��p��np��ex��d�J>�ܪ�HR3�PS�����Q��6���,��6-%KU_���l�)Lޱ��R�߉�~Dfvѽ�5�ϋ�d���-�L��>���U#��[3�̜G"��8QR���+e��Q�!��TѕL�K��3�LV�7�m�+��[@�/�����(�~O$xվטU�t�Ю/�W��$��RHj�8�%�Q�އ��G�y$u'^ځ��&K�e]�	��:W@�ѹc����r��1+`M	.�1�y�X�"��t��@�3��o@���!��*�Ԩ�>K�e��(�1�<�/Ek����{�+��
yv@���	&[Uf��%`�g���2�<Z��r��3,�8���͜7s�l�=��"+ ��1�8!II���D�g���G�a)9Q3�� 8����I� ��Hư�/ɬ�6w�}J���{���J��1v�\�̩s��'�������nP���(���M����H󖄺O�����0�Q_g_F9(���i�����`����Q���n9���yȴ�bY���ڈ��hC�wFb�!<r0�Qr��&7fSJz��KIN���]�2CXD����Z�9x���N�1j퀃��sU��G�A��8�%�r����{t,��s��3c�x(f�1�2��\�Y�]p�x�������'���s��!�&���v��U�f�؛��1�� ֜����9� 8�����>b��+&jn�����)�%��Tg����]�����$��ȼ�S֑�yN���-��٠�����[�'�&]s��mmR8`}Do������V��d���!E�l92/6��401ڍI(�d{n7�dT7+���Tb2Z�}Q,����c�XW��v:�fF�`Y,�%�|��~�u��E�������]��	`�l��r-19=�yf�	k���D`Jv�>#3
 ,ٝ����_��T��dGx_[mr��c%[,^�d��� �6�a�ʦ��,�{i=��}y!g؎������kG���O����6F��
�e�[b����7�i���Ϟ�G	a)ʎl��uZ��m��G��y��lU�PZiJ����d������>���-�(�����˹�(�>�@�8�V�{�u]���B��咋�\.X.l��)l���,._��;ަ�,nE�	����NZ�ϐ72��!� ׏�T�<��I�{����h򉝀&�M\&�$�K���J�_��ĉ�)��s�=ۭ� ��)�11*1����/Pk��]�eBԮՒ�u��ѽ�^�\�Uj�i���!3휱�<r��h�����Y�O|��s�0?ϴɅ�o?����������l&-�8��^ݻr>9j'�}~Ek��7�:��n�(�/����I�}l9���b��ޯ ^�K��5[�� ���6*�l\��ٹ^�����lfnz�����dG��h"�	#1��ʁy_���{�y��0=+%�ϿD�k��Q��i�����m����&�s���[ظ��i�zR+�:O���;#3�5F �� ����Q��L�<�8Jt�W�H�?:���/�X<#��!w��m���Y�M@oS -����b,�Ky$):?G�\��oN�����>����'� &@ٿ�+���陙����t<]og�
s�V$�0�ٝ��qq[֒u}>8�i�"Z�*�|y���-��c��:�����I	���*�w ����Ā���#��o�B��ҜU�&�}ep�h�)�&6m-v�0r@:J�cS�d�f��d;$��[�k�@_)G��h�:�O��HWR3��s���X�W��=��̓�?�S@囔ט�c��2:G۠R@O+�.�.�sF��jㆱ�Q��#�'��R4�2�&A"u�v��'рnOx�K[6f������>����}^�$��=����2�d���m���d2�M"5-V�ɗ2�T�������^��`q8g��կ h�h%?����-i'�!��2��㻈��촵S�W���<�mr�����;#��E�k�i�k��:�@��P�h)�2� � cJ�7.G��"�x���n���зʜI0�S�L��1��3�/V��2���O��������Ҫ$5�CJ�B�{�C�ߍ޹�Fo!�=㞵����G�L=#�@�L/��.7���&m枹ņ�E�2���H�~�K��w$sԀȖh�IM����r���	o�J_y�q�3�������x�������D��X��.�2�b]#L0�aKa$���n>���ÂI0��?9vDn�L�Ap�unA�i�����m��w����;��=3������'&�$syz���1��=��`�
ԡ�S�MK,M�𡟢��~�!8�e�������5�ͫ�(;�M\Z,��y�����w��RC�^\���xW���
f��q"�Ks�Q���bϒ��z`OB#Q+y|K�LbN�E��`��gEn�Z"�"mh����g{gƟ�G�)���*hb3��`x��W	OED���}�r������}����H�m����}Tb!1���mk��xdL��¯�������vB����j��|��9 ���`�hb}0�m�JiMl2���Գ
��`cD1��1�]�Iq��W4V
�`
	�q����^��W��4��]Z�2��4�U7�y��Uv��t��h�G����r�x�y9oD	L�~Ϣ�g6��D2�n�="ڂ>{ޙ}�ϟ?�#�i�C�k����2O,���3 �f��:���V�%��f��wT��`i%$�@sܦd�������ot��&ޓ� Yz�ocܒ�2.!F,�p�M�>x��ɺ�5��=Tz��5��-��-@L�,1��%�x�����͕~f��rzܘ�҄��y&]f��Y�lN���i����-��~BkBш�D1��rȚg�9�E�������C�)iRѾkgL�y���T��z��2�]��g {c��st&�7k�Ю�(���a]�H�{s�i��޵a-n���,��VmG�rM����b
[@F&8�r� �����&��<Ra�%����ahr�|1IZs�̳�رr����-�u�r�`Y\v�>����}2��H	e2�10&"F��Y�c�)������&8�`c*Ag�)����cɅ��[��jA�!J*k�a�B�Ѥ�߾�A��S�e;�[�	���|�ߓa-tX�
���Z�<d��YZS���s�?�5F5�SpOu�BDQ�r�!Y�ge�b��C�:���udҳR��϶���y��s�Lq�l��ӣ,��.o�����,��߽BZ����m���2��=3V�����&��͆1�
�G�.#\���qJ�&�$�H�1�@�����Z�"�["k�KW�t�z��ˍ���	�gD׳D�V��'	�ܘ!�*�1]��y��∐o�HlL��`��⮰�a��X>�E��{k���7��\}1 �#��/&����8,b�i�4om|���%Ou�c��7� o��%0̧�ɞ�h3���e���9��Bx����s�_���E�����.�՚�BUXpR�!��7��� ��Ae�ҡ���1+ٷ�9������1,�kʶ���ظ��V�^�����4沷i�Ϭg������̻��Ӗ�Z����l��������כ1����l���g�$��lZϣ�,L<��x�L��t�eq��C5�( �p������jlk���$t��� ��[�����&3�&��#J�u�J�Y�?}f-�KC��/&9]sZ;DD �Rct$U�1y�o��7&�l���ԧ�ϵ�f�x���=������HH.#N����?Z��٢��2i-
�tBB�U�t�;�(���ȣ&S�M����g1?���Y9�4������?QT�m*Y�y���{�=pi�x�H ���Ɨ���d�Z�èY^�s��#�RF)�d��m���C���~�lG�V~d�<s�h\�y'��|���������h|9��o-y��ђ�����I��Lyȴ6�kt��#RD��-��%��|H��l(fr �Z��	@�~ڑ�r?F��;�}��~��t�E�	���6���.#9�tF�PK!��l��2�������+H0��L�a�D2i�@@J�4���}��s��K�]����|r'�ډ�L��G͎�
O�#���]��aT�6�J�0:�g�Y�Z�h=���gd0�}=yx�#z?����8����wI�J�G��N`�M����L��lr!�@�\��!�s��y?z��Ќ��!�B����@��h���<�T�{���^��<}^Ov`S��o�Z�Vn���#R�&���t����Ƅ��T�q$3�$?K�oI��^~���4�����9����rA��5�!?`c�s���#��L3�l�����X�Al�7LzQ1,��s%�*�۲,y��`�"6+�l�7��i���06�ާ�k<9�5��>��j<�O���|�'KkG��[H�����N�ڷ����o�;o�i��J��E:�ky"i�X��&���Ք��cF�P*���-z�9�̎�ו�$� �L�GҚ�������W	�d����(���F}n,�e�71�?&D������6��y{�H�g���i����	�ɿ�$����wB������lN��q�?��fH��Qd8���H�e]f�$�d�������1F�n� R���X�=Jk��{I U���%�^�]�m����}j��.u�e����9�-7��\H�9Gc;FDx�����&��;bp˂�Kk����z� !�D<C����E��)'"�	��~�����º���$�'F� �����h�Q�G�@�V<~��1"��T��Su����1����V���w6��G�3�-�;���=[&��cn���k��uHB�;÷�C�KF�������篁EMz,����1�g��� <2���q����#��1i���_i�����eq�w��k��PV�8���'�A�����_�4u��-���WO�wcȴ��zC����9�unX�ɭ�J�ޓx<C��ϋ��4��?)H8�:��E&�Gk`�e��#>��{��>�?<]�g.GL;����`��bN�N�#��%X�IB�Y�J�).)�̥c�ǲ,i��-?_���7�F��Cc�i1!-�fv�gi�{r�a̺�P���"����8�a���G|h�%��\~vhF����X�>�|��.�3@Vat[�a~,�j��N��k����\��� =km���a_O�J�V �ڪ�����~��ԭ��{���1L(�xD(e/���4�7�帉6���uõ���Yrb~�d���L,����0�{�b����s����p�Xx���h� ������\nal����&�>X�`���q���XuFBܢ�5E%w1=����}�T�P�])��u�&\��W�]YJ�[��ղm��3?QyM�eI������������S�r@�럔B4e��h@R��3�)}����P@�.���G��#�8:��@@�S�%S����:n*��S�0Kw~�|�q���s�K �/�3�ष��iu�5��FV�G�J�u둹k�ٗ���v�Tz����>����8ʿ��[.S���� �:�,˂��Y��F�<�!�1� �g�} ��4�5X�W=�o���<�o�;���`�r�\ӿ���� ��)/������n����h�BLiJ�b3UB���;��nx��8�*ґ�ͤ!��S���(Y�Bk��ߐ�4w�pv�+��g��1f��j����lmZ�]o�3Ӧ&_XF�h=���Ў�E��[�^[$8q�A yL�����T���#��m����g�!�򤁽3T��g�O�M2Jf��/Ȕs���6��ť���Ҫ��vX�G��x������9,e{��n�O�xZ`���:#6�'K�@��)Eރ��{z�]�r�����9����	k-�����������T��R���!6�0�r��yÈ�eY�h�q�������MyAֺdF�Z �-��e&M��4��<t-�TۓG@��N�ޕS �c���"���<g���r�|V��x���ʈc��j����b����y޽M��,�c7��-���3���6#�s�`F�b0%���<sc�������瑱c��z-햱H�N1!ӱ1F��K �ת����K�Ι*9{Tj��Rw��fw�Z!�!% +ӭ���#}=�\�
�A;�$����I���x�ô����h�to�R[
C	�)��B��r�b=�{=�O��!��7QZ-N�������B2S���d`HL&=0�2# c� ��3�z�*o��Թ~tЧA���ڱ; �1�=x��,�5��m�����|��Z
+�&m���k�`+Y�(ƪjЯ��}�����rβ���)Sy̌h�r���1R���?�.ꂭ ���
��1ɜ��
���V>�g ��if<=�C����	��{�&�]$���C2�|�k��)�b�cP����������c�-%)�ʜY���B�5���R��&�SUfu��=�Y��>�?H4׋g��M-˄���~A�����Cs	��h�v�v:�3�������!�P�y�)�2�,�d�d�i�M�ǈ`"���D�_�(�#�x�{?��|V�盢��_1b]WX�v
KMe��T�5�f�K>����,H��d�t�c�g���sVj��Om��1�����w�o$X9z���)��5P��7�Α~��z.2z�L�Vy��θ�AK[f؜�q�n��Dn�Z3\?:�5G9{I��G���\_�2�Ge��b���%I������y�����T��3��'�|�\(�<E��i�
Ý�)i׋vG�t�5�>T� `�IH�*H�u�^���#�H����п�|��"� �\%(?ಓ͓1��T�'���u����{\�'(Oh�N�v��d���#HI�oJVf��d�6q
[�|'�����Ԯ���L!����1�|||t�w���Y��Bƚ����w�̝|X��e��鍿+�Д�x�xнɾ����J��+�R��3n����8K*���D�9�%-&��b�Ў��N[E���w1�F�@��c�e� ����c����O[Ȭ1���EZD|+��}��<�r�>F`�|���垳Α��6��C�:�Ţ#����2%�n�����y)����D&^�n_m"Ŋ��m]B�I6s��g�s)%8K���������u��!���J�����I��劘sZƐ0GƸ�YY_B���u���S5Ƥ\��9��<�@������R��V�sr� �hb�dh��lL�71��� ̗�:3��"���)L�S�@]J���v��lβ��;���o�)�m�2l@h�QS���v�#�-�GL7- �����BZL��,��7�}wi���2{�-i&�c��\{�i�c�R���C�gMq�Im���(�Hk�h?���@����hv��5w>���܀�>��<�
q�cnf\����:��(9�ꇈ��a���5 ]R����������`�����{��h'o�.g;��)� �����4S���jF���.�8�e�U���6^� Ji-ښ���*���$<Ҳ���<Hi��|�ofAX%��z�E�ԩ��7���I���10z^���>�qX�1SĚ�����f�M�#� �G���W���-�B��ц@nR4J���\��#���
I_m���`<�|+�X���%�y�Hֳ�f�k�Bx�c�"� �,���Հ��/�/��:*�������CΦ��e
���ϯ�ez=��;�m S�!�qˇ�v�#��"0Dꆡy(k���	E��S�L<�7��-�����x
���u�ծe ��KH&�3~�<0@*�����u�kVe�F����`�~<r3���
9�����Wc�g���Rm��3�~�K:�ᖥZz�(�=>������G- ϼ�g�$g$�o��g %��֎#�1���Ex?��A��z�L-z����&��u���k�sz�T��~_q����_WDXs��Y���KY/_�d��+�m ��3�D��ѣ$%Bȿ�P"�����l�0p��1�&�4L���,��w��\���r���&C`=���2�#���^)���v�^�=i)5�Z�z���5ŗ&p}}��M�}k�����f*WT<�T�}K"����mzcD�sd�������w�|d���[������=l�@���k͟�|]���g��Y��e���"�k=һ�/t��jה��tO��r����w��o��2:}�Jӱ��yEmI���,�����-^˼'# KyD�o|-��k�e��8��/f�g �6xĽ|ΡWz@i�)0�,H|�PII�;�����Aw�ь�@L���[m������ή�-$�?n�9�9Vc��\.)�,�2/�z�/�7�L-Ld�
&Q�Wn�.1"X�BA(�Z��ͣCK�Ps��|b��uRBX����#�H2���B�_N�ND���>-�l�����]�#��`��lD��b��W1����?�Pj�&Z�����m1�'���T9�J+7����z@�;�,�%=���A0�~�5-�|F���_�	����ϔ���D.�w�<_f�z�f�lI��\5�:S��N{��「3�?JPN.B�pr����ù-����~���?�ŀ�@7��nk�sTz�����m 3�8)��<�cGc�v��0��Q{G�OIU�V�|�r��	zt@iɉ1clŜ ma�DR.�4�u�ȅF�ӣ"L�9��ԥ��Ŋa�)��3e�f����&�ן���@_�_%S�ه��{���9��W�q�vF��l�x���!`R �tI`�nM����}�TI���
f� �i�0�9�W+�Y͉�>[��_#�c�W-o�twj!q�"ƭ�Ve��P�	2��=��v�Y�]n2�c���#A��JC&�m����c��9Gc�@���X��� J
l��FJN3G� nR|v�΅qk�N��t^���?�*�����X�V���Ö��#@�H��;w����B�#[l�(��w��l�h)�v����G��3�
i6fK���~|�H6z��z�Re{�YT�S��Z�q�'9e_fe�,�>��N���z��F���1\�:�"e�����zCm�ڞ�v=Z�U�}ϼ����kX�Vg�����51gTi�!���/�>����� ���������l��V�<n	ۣɃi��ȃ>�����5�Ĵ�r�����傏�����4՝�������W�o�f�A�x+�0?^��;nV1JE"�̏&M���M���hY����'�bs}{���(�ET[<di:�$YK@���x`�L��Qg�cg
��@������v>)jn��v��3�dh"ۘa	Z����[��W��m�z@Q~�׵9���=��g.n�C��Nl4�=����}�8~_��g�=g^s���d/=˙����c`f^���~�������L�-�C��/�~�e��w���3nc ���˽�M��N֣?�Ovm�u�|}i�W$�HO%���6� p�^q�^����*����G0���X\r7KTW�S�L ��x0������G�x�1���.��N��@�\�_�@LA5f5�({��d~���AKR&H��������O�̮��:���Ή/,ԿGA oG��~�-��J�+w�3`��>��1�"���0�R���f&MZ��/�|,p���Q�f$#@؛kr?bZ�Pخ֜ ��F�~�N��h�~5˹>An��Xk�l��K��e�|�J��]�9H�����{��oK�Y{������ �J)U�F�i��%��,�h�j������\�D��v5�S���q}Bz3�8��ܚ������fmr~L�'ka�,���>U��ט�\a���Sn&�`;�^�Z���k~W>�.Svʓ�P}��T��2j���w$M�P�=+��+&W@�=gɨ�#S�,S���f�u�P�G �H���R����^������w9�]7��/��)7;�q�D[�[כ�g7)�6�Y x4�{ �'����d���فI=�X��}��f@��r��/7^�]hj��E��c��%������?�����<�<����8�����G�I���1��?(�o���^8�
W��H�TV
��"�^o3��������/d��b@�,�S�(AG]҄N��6&0JIO�Yv��GC�5S�u.��qaoV�B�_k���3LM��g;V���� �v��l��%u��$Z�NM^�)%W�<J�W�ɇP�����]-8 ���E����E�%g���2��L�3m�Si~���Co~��gD���%���3�{���D��.:[�W�<*��O�|�w���}ɱ����E�S��*���K�VA�V��^K�f���p����z��F�:�X��ڭW0b*{�1GEnZV>�x��WnĎ
���fU���M�3y�O�X�͎���1�1$J�Ԏ6
�3�&��~�ӾX����X�[X�@�?"����B�}��<�=���%D���G�>�-��1� � ̬�k�v��^gq8`�&�����h�fc�~ȝ��l�#�)�n��U�#����v&�ܺ:Շ*�^H�%֤:����|�Mfz�����RF�N~~T���-���"����'�.�����"YMjG{��%�3��i��Ŝ[�w�[۰�qF�l��!`&�p��X1U!|~~�|�t�#��9��9&����G�r�9�G~�t�����M����Q_X�S������d*[zUӕ�jG��~�9�wK����$}D,��t�����97dW�ߧ��azw��1֒��Q��b��Ǹ��D�zG�1rJs;}q6�O�=�&��K:�t�Kֻ\��\����&3�Ȓ"�S��� ��L��p���4�k�O�0���"@������ْ�����ڭ ������,
t�4{J�6�n�:<�`5�B��Q;��|����]�\O>�^ۜ!�P��{�Y~�c���;������˾i}����q��7v��k�ڒ:���J�����y0C":8��YTM6��^HOmy.��Qn
B�S&�Vqi	���^�+-9�;f�lTۄ���v�g�%�n�?E�]^̘~LT1Se	��{LA0&-���4�A��Ci����'ų/�QkG,���d�G��uf�����O��� ?���r���tȺ��'�9;�JgdV���������}���}�k_�O ��͏�w�#���\$�j͑�s�߿r#(��1�����ǒh�\��6%#wD��H�������0����*8�n	��g�x���\/I������c�scl����>�5��.��v@�W��hk�t��)#R%�T�<��%bJH�S��kk>g\�5�:8�3��>WA��+��} 3n?���If�t,=���{�_f{����|LQ�!BZ�f�Rğ<��Z�8{����Y92g�1��y��L^1�b:?����_�19��$�3k?2�4F���X��u]q�^�l]Gu�P
�:"��7��N]����Y�R[��f'��9(ƾܳ@s���;��i%ɗU�z>��:g�g�)k*]�b)%[�?�։�S�\ā��$<5/	�E)�-pq"�t|͹q4kڞi���k�d˹�����J�{zD��K"�~�1F��Sۼ+)�h�~'y�OfB�%�i�҆��2{IҘH��r'��Jʤ�̜ƺj7@�Y�-L"��C��#�J`��J�0:����#�mQkU���i�0-�����oɿ��V�H������g�g�i�i�l�����gN�([�����6�T���!�OIϰ8WX@��%�#�|����܇�z&N�_�U��ֹ�ߣ��d^�}�z��uF�\|4&Mk���=�\+�)et����#F\��3* ��~��
`#ۋ���)��<V�W��ef,s�f���X~]ن�GM�(%2����-!iCdwUzZ�K�TtfH�L_pFS��{���Ki4�������gKz����d�ec�[�z@�5_�����{}�LL�=�N@3"�����vK��5|9C��w�s7!�@���M�� !vԼC���H����$&��$������؜�����.ay�Gs�5��^.��y��M�o o.ۑtB��`��� �v�)M`�JV�@��X	(���
�,(R���ڪI���G`��i��������<s~��is_�Q{���^��h����H�5+�G�[d�M�ώ�d��Nc��\6L��l��(�׸5'ƀkwn�}��tv3ut�z�%a��z��X��Oc^�q�3�c9��9[��[ޘ��#�������=g�������1���l�<3(Ǧˌ(����8�p�X�S�����s���2E5jm�[�!�`5�1�ܐ����/S�����e�'�~�B������ؙP���=ʼ�F��2��3R�����=������8�\_��zD$ ��޳@s�]�TeFe<������g]Gꀞ�<�3��)����~lsj;�t!�Gͦ3�ǳ�mTի��������{ϓ�]��<t.��Yka3�c,\���Y�m���re�)�Z�@����>�x'����Ǩ�XP%{M�O�I��Y.>�#hq=8��n��ٴ�}F�V�%L�L5��6p���>�rڵ��U�^���b%g��gr̗�D�c3zY��%�$�!������L0΀&�Vά1�߳2��uyZk-~��wX�`l�=+����@}f�:�֓�f��R���_̲'�N�����<�g�f�#>���1��G�̸��� �����5)nF9��,��lm�4�6�Q�V`���UY���n�{k&���!Wչ1���7��[>��&�3���v�#�b0��G2�pc:'Y��rA��4� ��:���6�{��-�(Ɲ)�-ۣ����ʎ�(� +L;-�����fu�O�W���u�}A%�:�j�@Y����I�7��\�&���d����{�88��|�n�Z��r�_W���y�e'��K�lL܃�_��dd��1#�4b�9�{D�m�c7���"����v��-�4?S���l��S�n^e�6~��U$o6�AU�`�.��&��W���@���#`�1w���Y�%��p����Y�70���bzQ�s]�|���~�iٺ�W�q�G�{���&��W�M��2���������u���O�D��$o��L&��bD~�l����� �Y�9�`aA/
�!""�����+�bl�F��P-t�(~�+��3)�_k"M�L_Z��3�yn�����"%߻a�J��/؍�+���#��i^��ǳ�*��P�-P�6���=��ߊͩugcg��R2F�3�ԇ�W���R��%�«,�p��7Y�z���YL��R�J�ԣ���XSW0r��7��1ycsbL,e�ɌHTf49Y{~��+`����R���)��]ԝe���9�X�׼��N�%� �Q5���GPRg�1�)�������l�������MO��jcK�$��L���}�Z�k�,�K���J^=ʽM磛�[fޟ���E���,��f6\�j)�n�g�c?6[�B��=!�Q��p����u{���w��n-��n���7���y�6֜gs�kLLg�:��\q���|���V��)eKz�Ō�fy��=<��s.e8�n-,b�-zjgM��z��n����*&��k����_�g��T�x0qvc6���_�;���Y	���\T�1�6<2P�s�7��2i�~�����7�)���߹�ĸ�5�y6�y;2e�tn+�A{~��g0���	b�	�U���~�Hi��\I���ΉK�B��&����#D�c�X�����L�;R��,N�q ğ�H(��WY��J�̵�x�A��B:F(�!)�v����p�ͺ�a�����}�]�C��'!�'3��a��l�9� f�ؔ�k���1,! 80E@;����ĘsSE�b�HK@,M�絈b����*�S�A��h��Q?�)~Vf ���9-H�(��$s�I�ٺ���/��p�DV�߃�%!u���i�6bln~JАbb9�x�4P����9��1+�\������w��cJ�C�^YDb]�ff��]�����߷6�ڽ��������V�.o�C�U���M Ls���,{�&���V�4��U|'Ct�A[/@OS�eI5`�۴S|%g��o>�Y�a�^Ɍ�������V��c���s�swz�Y!Թ��?<��:��M�#(��X]�G�����~�a�������B�[�u��"έE0��.p�߲\S�K �O��o�{Ų$���l-kߋ�~ȼ��R�i�� ��M�6��bb�Ʉ]��h�?�-�߯�F8�u�G��]>�������?=|/!���ʿ�E�vr��g���g��$��ˎ���I�oVJ$�Tk��#%%{��w�}�	xx�)�����R��Ƌ�vLQ�y�}8�\� �$@�1q�r��YK�����v+�Ʉ��L�P?�r_!f����h����SZ'S�]��+���0�����L;�?�2�㤅��g���ԅ�EZ�uO��X'�T�9�������c]W�n7|~~�~�]��g��	a{fe^ c���}���>���(�+J.��1Hd�R�+���z�6�<ĜS0��`���Q�D��h�B�����%kQ�����{h>*|�7bN��W�L�*�8#1�-��� $cL�LF�aZ��kc7��r�t�z��8s��q��8�Փ����ʪM�>pKcjϜ?�� ��@�C�'����Y:~,�[7�	��k�}�\R�}O7�{eQ-�Z������o�-h`Z��xղ?�o&g����Ii%��C��Y�@�k]W��n$2�"ʂ��|����J���s���t]�.�>sy�e�P���Fn����u�����5����Ћu���pnY�|\��Ǐ򏒢�v�#��"n� {q�3�i�hZ$2H��	�S��UneQT7YT���4i�x�L���fގ���l�.�$t�m&Hf���R${)�r�N�g>��bA=iA��K��24�;�9;
6�{��4M�\|xYGcL�W�zV�x�ޣ��G�OkLe��2���ۙ��D��mG������-=eQ�}rH�n@s;n̈�u#]?�)M��\���ύD���J�N���\sn��d���5t�A?��%����m Ӈ�C�x�L���'2���d�^>�o+.�!�k������������kj*O�gͤ�|6���W\?��� ��&��2�e��-~|�k-^�;`so�vvI��3
���֖D����V*v�'N�WC�����9�~�33��N߄U�`�̩�:�ǒ�@��:P�Rp�,&��<�ߏ&-���{��=�H�=R�L���2�3�#���%K���� M`����^��'�2�������h��𶩝-f��y���,�w��:�ݑ������������}�l"w)��"7��5��E>����5gE�AZL�Ǎ<W��R�#�y��Kψ���':nqN�=H9~�����u�����Uם�~��~.!x����� L�˲T���
ʓI>䔾(�XX���C�����5����S��d ��L	j�DP)m���,�V(`�B�1�b�p�g-����S��8�<*�1�|n���C� ͖�~V��s�^�]]xS+{�?�|�WZ����F�/=S��Rm�+i��<�)��l2�gA�ݑ��Ys3q+���!������Q���[.�����Wy�6���U�4
Hl������G�Ah��1��풒�����w���ӻ�<��ov��J����Ioc�]���k�7�d��Ǚ@����7?���O$L�	�Ϻ����a�f���`�]M�� oMaT�6�g����De�A�'��1"3Q�;��H����`Q�U}�
���?��Bmk&D�\�Z,��(h��I[��	���.�� �J}!&+��OlƧ��!桗Ze$<�l[�G�5��zLj2턪ܦ&e��"�K	��=�ȅ�y�'}Z{� Φӏ�5��4��w6�ӣ"�EI���(`)�}.�ԣ9fi�ɣ�w���֔���mCY0xz3�2s�(�NM�X�I������a�����Μi}�{�� l�Z�V�v��ٴݏs�� �׎���E�E�*pg�[��@�"���@	�	x2s�LTZ�9;�\~]�MW�6�[����sڗ�r6����6�F�(�#E�@f̋�X���vL�j�_�a欖��H+K*M� ��'����c�����`mv�D�nԼ8g�mm>x�SY�Am&�%g�rqn�@�]һ�6y�ki���w�|�EY3��8��$n��s?�)� =j����))S�h��4�x��WJ�Odp����ό�<���Pj���7�v�m�[�sfS���-=�Y�AZ�v�(���g����[G�r�k��IK��&f���b�B-໥/�	2r��H��rU����q�Ѱ����"��� ���1���\ ה��9��� Q��.�`#�L�|��&�	X�ha���!��ˠ�`0`����/����"?��3���GǶ��3��J�	W��B�l�<�b�R0�>�f��+f{?��a�'.V-� _]cg>R��O�z�����������a���L�<����R��;��E�r��q��zӣ�m[�L��}�\�j���<g�t}Yň�����M�y?����s>�,�y҆�'v��Rr�8%_�N�`���/7D�xi���V�^���̦���9e�k����y���� �mim������d7
˘M����6>���9n��|�Z������L�P�#O��{��)�����yIHc����`�'r��T��,��Z�%���j���0'׭α�Х10��0�X������cv���4�k���֦An���<�[>3t���ґ���� ̙~�X��s��7_KJ��bh[Ɉy �0BSQ#�vV
��o�n�k�[k�-R,g!��3D��g�N*~P�rH}�9�a�s- 0s-n6vʵ[s��}�=�y�H^�m4eZI�{�ɿ)8b��r����TbtN�}�ͅ��sN��eOm�+��ue�ǅ��|S��E����v6AZ	�����R>��lO�Dy|�l��K)��<�
	<��|���N$F�6��f��4qZLlnCJ��w���̐*�T�Ġf2�A4(�z��%�&��P���D;���8�b�����G�Hő�o �%ŴnmQf��x���?Z\蘒�g@���p����%��m�@��(3C����Ͼ�B��R���%�:�e����>�$[�L�з̢�w'���>�e�����D�Jߓ2�cl.T�U�����<ΤJ���o�L��9�g�{)|4v���,8`�mĸ:Y>x_�q�̤��:?�H�#	}'�9Kx[�G>}W���?���K~,m.��W��3|G7]-��%7�G���F�<,����G�!��� .��}�>��t�n	���dRl��N��4hl��C����wND��A;W�1��~W�UHi��ͣ>J��
�@���̄�J��9����<m�4��Q3o��9���O,�^J��xjf�#AF21�Yle���j��,��Nl^��r�����Ƙ�fiF$����9��7��|�Xi~���l鈸���硙�{}��n~��B�}��i�՟�vK��5�W�-�n�s����>yb��r����6�N���_G�<f,�|�=?�I�<5��N��� L@����x!FD���e�{��,�1���l�[�̣��8Ɯ9'n�fd���.XB��T��Z���
�i�7�Jv���@��58�u[����v&�m�8cb�X}(�-#����]ً�&�T��oJl�`Pژ�nbV�t/ʱ>���ᖥ(�^��H��jm`Wr�)���XZ�ii^��_~�h��3���_��b�5xK�!�ی� ~��Q�F�0c����J�	�<wm�1
�qp�4io��7���(���M�T�P�"��5n������ׄ���Ǚ��S�ÝY6�ҧr-�#i���e�r_�cF�`�����\#�$Y��/���coe̤��T��gƖ>��|J�����~���V�ת�����m<�|���M^T4��ڬ�L���(�����1
��1�m"�/�+��pΌ=~_�\D���Lί�מ��q��q���$�dĿ����,�-��WI����gun�����_U���<�y;��{bBLlք��W�Se��Ш�w.Y���y���+~�d���Y�~�ίZ�buAa;�m�����ٿ���w��&�H�Ȏ�%ń=�����Ĳ�,�;���ڎq[����K�m�n����C�x�R;��x��|K����T�h,WI2gm�z`��G[1�G�Xsc��;��=
�/�V�c�d�䖙�%2�����?tn�:tm���u{�꿓�)]�]��6L�|��猘?%���:������ؗڗ��ɸ�JoC�?o�/��5���	�<6>�Xh���E�&�M�3cO�!Ƒ\L�����?*f]�=Wi���F�5��~��3�%ۤ��dP��6n�@���c~L����"�f2	xc2M��eq%xg�����>��l&�ݘd����� �s)9�щB@��~��JM(c,��w�g&g�C�(m��^�oU
���[�ֆ�����v�9���܇uݢ0�ME<�S�%LmCXy
��ɬ3��r3�f
*L��8�Y��+��;�.J>@��G�� vF��#gji�|65p��/7\�.ܴ_6!�;�S:��9�le~�Cw�Ƙ��)	��i�!��I��B>�lʼ���svn���̂8i�xք;+҇\��y������F\_��{e{z�U��O>#d]����҇@����P���Jk�L?ʽ5�g~��oe�>�#!�&a���)����mXk i� �Ol�! ��`M�Y���KI
$+�|g�� G'�������dD����󔠐V��K��J��&��K��<gDѧ��W���]�/*-��U��@3���׋�6�co����&Da���q�V����m3���{||�:��Y`�jb����<x9���
���6Q0�����}*%���$S.�@���L�zR ��tp�o��`��f��a,5��m*����T�٤^S7�/gX{�;����nS�-1x�7)�M�z6~~���V,���Xh4s,m��2���m��67}��7��@+>	ܭyS�>w�V��_C�ϵ� ��j���7ц^��#S����\6hxO�̹Aq�
1�Ǹ�&�fZ��W+�ݷ�6Gyk2��{�Y� ��\ɿҕģ&�8m('�v���^�A9��.�\�dg��4�G�1Ҡ\��	i�l���{�R��_w�=i�u�%�i!�C3����-4�wb*[�)�g��-pǣйW˴Mm�b����O�AM�)��;�/%���H���+h�,�����vc���O�铛 �"��)٪��	���'�	�Ɓu��4 �q߹��M�=�Ei��J+��
zc ��
hT��i�%5:�������g�9�d g�e�1U�/gd%��2��<���gb�n[�l�FU��Y�Ë��H�-m魑�w���i Sn��x��w��α��+�xa��s��d�]S�^n7����?In�[960�Ǵ���.�|$}�WX�"���qY����+��06��c"b\��G�+B� ���Bx��Tu�0��)o��N���(��V`�l&�>J��E�h�1�wzi�f6��uX���:CV�ʳ�wt��<Q�Daj;�cJ�� ���:�T�Z���L����~��f�Q[<��#i"Z�	��;�?�f�Vl�+�cU&�G��� �־Liq��]>B�����Qؚh,���&-�E��Vd��2��cZ��	�M��u���/E�4?ˎ@�C�����F��'�!�2���rV���g���V�wJ߶M6	��V`O.>�	z={�҂�u��-��q�ݦ�
�VI��v����a�-_���!��2���)@�$��+�L�� �����bzh4��N���	(&��5;��GJ2T��df�1��3����܍nY���>P��\�H��h�T2���GE2�e3�(˲�u��`�re�f�3zڵ[J�'��,�� 6aRԘp����l�5�wՍ2��E��+���#��=�ڬ�gDd�8j�̷���xo%{o��ք��6�U�o�d0Ne�{���V�ٙ7�Z �b"L׬�8�)<��v?�2
|j][�2Й��z���#f��6��򶟽����!zdIk|��O>�v����|e����J�tc�,�����H+�Kݯ@������o���5��`&7)�䩔R �P��j�ڵ�r|u��M~����;����?�ۡ��$*;(��r��c��ux���=}	���<�t��Y�h������Ui �o����ے�'�e��R���1����>t�/�|ϯ��7��#ɫ�<�$/��?"�.}%{�&�$��یwF��]������m�Rj?3�8��~�H֕����V�ՏH+���d�x�̆1+��yTG0���qK ��hF�}�7Y#�}��x�z�.�N�$�ש�o�*��Ġ�X�����Yk��J)�zy���^{�JQk��ܳ��#c$�6���>�Iʍ�O����YQǘ�IR �	�B�Ƙ�d:� ں�Es�i<��lNaה���C�J4, ��T&��_L'&�d�f�̖���?�?$��������A(ݯ�6Je�˹�l
���\�U�.g45f��n˔M K�n�>��'�����1Os@���Z߲bN�.'Z�G~m<QNA����u��6o5`�b��������xT6=��' ����|��>�s��>���D�%+��I���y2�z������Ԣ�c��g�j�UN"H�v9.��ڲa�)��,�t'�W��D�0����$����-��{n���r�_�*J)�Hܲ���1nI�cD�bx���b�ό7��?:m&�{�J��#|N�uf��3� 3�(;��iLJ5��N!�`���<O,&Ee�U&��r���E�<UǜGZ��b�= �5V�hV*����Vq���
!T��c�kka?�G�����Z��G��~���I�iQ��3)I���J�5b�4Py>�3H������G�
aȒAC �K��!�9��=�0�T���w��`V�o-��z�~�ʇo~)I���ۑ��Aդu���tO���t-��-H���~j�@=�����3�ԝz?�i9l�{t�ү��yf.iM�ۺL�ټo�����1/�k����β��Q�hb1����.��,p��j���iL]u�9W����D�����g���G��L�+�����hx�1��o
1��Au�^��㾒$<��1��k�R �͚m_K��/S`�Y�����M��Sd��R?�5[�l����e2�ڻ��U�, ��q%K�H����-�8�_k֓Q�ʌHv��>�G��^�Yj�*�Cc�x�}�� t�X�Y�Ǔ{ 6�	f>��"��߷���lS��Ԯwda��*��=oaɁzo�ݘ��L.�ܽGEZ��:ҿf�g;��$�Y�gVcv=j���Ϗ��#]�����;��H�~)�/�u�cm�l��b]�3��mv�~YS%���ފ?�H�%��2�a�n�\e	`����v�%���?����G��Z��j֯5�Z�H����af�k�-'~i�s�y�*8�vDf��f���yF���5�K��,&�G��`n}{�C���L���3�ͧ�vYvQ��(|�2b�ZQ�t��1TL���rd�U����'�h��r7�kʾ�����&��I\���ˆ��Ish�-��������Z�As v��R3�̙3欌3dl�������lc/�˘Ժ�5B��|C���L��ge��8�`|Ƭ��]����k2����|~(f>���1����<��v9{G&���@ � ��k�@�H�u, -LL�� X�0�c�"..E�Z,Kr���  �X�hM:_�MHy�2�p�^��ǆ�&w�?]iH� ��]�ym|9�[)�4��^��$j����M�Z���9iI�Rb_W�T��w�1g+p��t�V/�r+y��ç���;����:"h��z�]}��e�6��-% f�����QVtl�
��������$�/�Y�Z�P���s�1������' �����=�}Hf0��zl�\'�AG츑TANL��˜�K���yiLɚ�@`�1˥E��M�(���EZ'���\$ �B�Z���5�[�Ec����+:������,d��|��؛�t��)o��͗�#��?����ǏR!�w��~����CҔae�s�^˹���_'�<�^/?p�\������	���{_%o���:��1���30����b)9�X.���:���&o���¾�W9*R)jl�3��y�Uy�_ψ�������>{E9���_�R�rQ����W�k�~9ș5u~�H�*}� 2�*�m���DcD�㈹>���le.��V	R�j�|Ue�|�}�ş�rjht�wg�B��:s&��Zo����܎�kAP׈3E�fcL�ԓ���Lʵ	�7ǁc��Ge4�ӽ�M�b�`��A����q�fV�uM`]�@$�������8��܀�s^%��� M?�0(�?�n�ɑ�q"j��&����2F�<2��R�A.JBv�Rb��{f�<UPX�i��_�\��x{~}`�
��W-Fg���w�
Xi�<��v�g�(����r�>cu���\	�# e\��1F,�R��K��5�^����l#]��\��B~�j9q�HOB.����=�"eϞ�_i�d��t�<kF��.��v2�����>�;s�9��zM��ۖ��I�8����^M�%LJ9�(ᆥaa�d���Ԯ]�"Ĉ�r�����_���#���j�_-o���9�XS5GČ�s�r�S!��5�xV�u�5�$nWK��d{i�m��P�i݃���k�M=u�5�����V�Of@��Wt��r9��U����G�J�r�/-_6i��_g�"�a��h�����~���3R�{�Pю�{ ��8礬���'��m,l����$�=�LR�V@strC!��W��Y),kL F���ƪ�t��Wmk�B�W�R�I�ַ�+?�Q�z���Z��K�i����rm���{8�uˏ]��N���I0�w���P�B�!x��q��q�������?��_�����<'�+��-&҈<��c)���X.��/ ��r���	��e��[���Yü�v)4��s�\. 3=IU{�����L��`�Sx�;E�;2�ӱ�j-є7��(�?~_�}�X]���ߜ�*�3-��*�ݻU@��?�y�(���R:���e`S��] ���"����f�d�x4�9�1�����c�ș���2�D�!���C{f�lR��aKZQ��O�+�/�|J���g�g|,{��Kc�w̓��!��gkao�k-��l���9"�vt_��_��b∌( &�\M�Ē-%���.�:!�[�z�knc�$J}���l�ķ������K�N�W�qǼ��dݑ��!�*ȷ���w�88,�aY|||�\R��_�w|~~����q�����/����3��W��@&��|��k5(���0�K6c�'H���<|�!��H�C�u7�'��Z���ɼ,Ģ�^ĖY�xtDYi�}ob�3���/��,��;�"�50�*=*�m��	E�WJ���9dX*���7j�����o�6�- ��Hi�Y���K9w�@�Y�<pi��yK�R��R:U�K�̲iqe�҅����u-��#,ج��~m 3x�ˠ`�f%�5eks^�:2��ˏ�z�w{�y�]H�iΥ���(os�mL��/�c��n𰉭��J9lc@����"�a�?������<K��I?�i�ߑ�e 6�L��)��wq��E�mU0x~L8�6C�@��WILJ���Q�t����'�{��w7R�y;�x 6N�w]�l^ۢ��[ kf xj&`l��|��fLb����vc_˼{~����Am�)��v����q>�8O��N�"�������ا�?h��M�(�����T�ZOq�Y]?�y$ϼg@�y�I�.u�^�>jr��|���/�%�(��m�����#L�0H������0��e�������e}9*�Kads-j��������`P�;g�I*���o�\3���^ޅ8�`T���P�~��-���4��������"��V.*�������F�.�f
��43yU�6��#��a��2��ǋM�����]�d�����g����,&E�3�<�4%U�g�=�P�=hm�c�����������˷�"��}�'橩���~�{���!��,%�#�O�T.ay��ۅ�[��P-X>LZ9`��>?�Σ��Z��o=��z�f���G�2I�����*�!P�GZ`w�O{66���cs�gs(���ʜ� )iK������ky=>���#��;���S��������޻�!!����Yq6��fq����&��;>����[o�m�Z�蓙ee� �r{A9O�������l��vF�
l�=��^�s.�+9_��z�/.�9S�VR��)�� 
��ŕ���ౄ�l�E���i�����j�d��foUP陥5�*DH!��;Y���R-Ty�;Ȗ�MȾ��5��)��G�苮���Q�1�}���}�6�}᳤0��r��\we\X�-�7��y;��@�&Z�v9Ż��r��O�lfٚ��mAx��6�#�3�ڢv�}�;̭��]���???��s�j ��������0ϯ�@"�\b���5f~N�$�BwV�>En˞�����Б-��)�������4�6�۳"ǈ��+w)�\���ϧ�v�s;#�(�'p�k�4�/�hJ�~��W�Y#B�ekbm����,x��Z�e��Z��^�^�@2�ǐ����l�9@�'��w�eA��}��Nm��Y/����0������uXo7�����N�Z:I�XVr3��"cbK�u��"��z�����Tv� �0���!T����]R��eYp�,�O)�h�"Q�6%d�-�|qخW+HmѦ*)%�K�L��960�ڔ&H2�`���)�wʣ���,@�A��9�wjt% ��R;�P7��Sp��� <𓾘�s��j#��� ��������
+�*j2�G���.��O�ِ�{�Y��Na���y� �rM%�m�FGw�SG�F����=r����曔�˺s�\_+�ɟc,�%p�!V�þ��Ť�Ea��j�g�����u�K�"7"�3[1Įx)aR�������)o���)���i�L��#�Ӯfԓ�Z�-�~�>���naw|��,�PJ6%ߕ�o&�&!9���i����=�̙�'w���W�X��3m�v�#yw�W�lpN���Θ�e
�V�b�xҙ^c7�bD�+��¤�~1�P��mf����1����#9�/M�R?�V����������b�W���i=p���&�ғ)�#��s�j�6s�����ti�WR�L{�d^1���uf%�ͪX���8��_5��K�"\ƈ����6����a�������l�@G�Ɔ'��ϖoUI���H"r�*�L�F���ǲ�H���:ɎXa�y������'~��	�\��L?���iK�Jb������>�H�n�ڕ����(��R����N�vL1��>"���+
�sK9������Rv�>�G�b�[5��Ll-��(�R+�Q+*���H�w_�*�徕��Q��V��>�';��,��gR�6�[:p�-�{��e��[������}�<�=��w��l|�{P��e��/�>�n���3F�|7��tW��}l=_)҄��[K����H�����Ac��Mc�`O�=y])�\#B����y�X_-f�Y���'�l�3�y��52t�A"�l�'��}����+�� ��
-"���
N�&���7HDsژ���=�R�&��wXk����p��~_+%���J{�:��9�����YTO�}�b�U�ނJ�29�+S�0��EJ13���v��)���M>�[���	l
�G�����Q�?��G�|������?�P�%� �A��I���b1ez-~,�D��:�kn~x��-�ϫe�<\1�@e��ƕ�����j$6o+�C���9�̙���-�<Y�>'Q�.�;���K�y�<����'���-���M����M�\:v�B�A�?�ͱ�S�[�����s�<���!m�|=@4���5ׁZ�4W��탁��*j�,��Z>O뮯�+��,�g�]�Z�5���X���y>�����ǚ��e���y�p̧�:��͕i�c�(��-���`���G��������e�caږ� ,9?�5��m ��ϱῸ�B~љV�-�i�)@�7�R�$j��*Ҥq� �Q�I�ʄ����䎑�C�w���&(-V�?#'�9�u�H�J��^��ػN�i�#�u��WI��67	�_�2y?*�$��������Ȝ�`���1#͚G�C�bcLY�ɹMD�fg��ݯLe��-�+ѿz~؀���7���\6�~�8c>�$5�����X� �G������[Θ���uv��~_�g�G�o�E��^��^`���67%��h��g���^P��{S .�W�N�:[R���ݚ�@��{Dk���¯c����Xr���R���S�<��������4@���^5�JJ�J	O�	� )W)	(��}�wEy�F�(S:���%F�m�w��,����ͳ�H\!p&�����	}G����ڧ�F�b��[;s��}�{&>�|�y���m�`��B�&��P{-_;e��I��Y��H����3���������fr.�y.S5q�V�K%������\�S�FWn����rPI���n���3˂�}�ɴyFNR`�1��6����𲋏�
�N��s�1�̑�}�K�����+_'�h��pp���~�֓^Ж�x��V��Qg,�}�k�3�6���+>���c�n���	1���9O�C�R9rq�Ќ��|sy�
|l��@h����Ğ�,�m���|B"n����vp.�w(����֓Y3���?�݊1V�+�`rd��xi� �iI1q7�Ib�aS$#S�|f��M��az�bG̃l[2�:Hޛ�8#������>�KR�ȁ"t�v�S���=�~��k��y������J��zԺ �м/�{|�T,<�w�T-�d۩��H*��;��,��5=�!>r�!�=����yJ��@^��V��A��d5�S�XK8[J	ә���0��Db~5yt��ѕ��$�'�{���j��d�"	�G�2�ІǇ�R�a����T��W���=c�M�T��vք ������sXr�ǲ��Pn�]�
Lb>��}����5��Jx�5c�y#��TJD-`|
ipX,`�G�>�}34�B	v ��/ D ������Ǐ-�1���ZL�֚b��ٴ���k-.�Kņ&E��D[�-t5�eL�b�����{�g�t��3-h�~�*׼^/|��i�I�ߩc��#!�#$�gM���n:@�5Ak ��9L
o[�7ET�p�����͞<�F%�2����;�5E�s�P���9�F���i]���@L/-�02��ܖ{��3������P�"ҵ����dU�VZ%~�_|㦁#v��u�o1ox��� f9�}G�;|<�>(���Lڌ�M0K��ɇ��E�����R#Ao�ؾ�]��|��zdև���,�1�J#��&��aIo�Q׾�YTx{ ����m�1j+�������$�\5L�3,7IG�\M��ܧL��84 �!���cM9�c.�RKD�,L��~�����:�3fH��ޱ��JOr�S�K��-��Z�����۟�������zŏ?����~����߰~�2^Y�2E�,ĸ���CFR��{xc&|H��!���&�6��?..'�unI��fA:��#�=�c��lal����K���K�)6@-�gxM�i����3}���ķԝc��+*hM0-3f�����-��|���}Ӕ�ȍbTM�2Z����*�hc��/?K����.[�c6߻�L�Mb�Nl����6��=󻠛��:�ǃy�ʣ�M����ul�Mb�}I�������a?���!-���P�<�RsD�0�J}�b75s�֟�m*�P�u��r���U��[?��
3�=b��!B���L�<7.	�zl�c���O�&�5&���v��v��j���o�����~C�m���r�ik��ƑB����|UKG��$���PYIl$��D��9�hO,���)�ƈ�.�QE���h��+�IX���(�Jm���̃��}�%���9�)o�3$�bX�{���0�J�'���H��:S�?$���A=���6E[��1py�?R.L҇�� ܗ��A�8���a�� �٫t��վ'�}�X�I׏W���쌍)���j��~�327\ǵ��ʣ���(��,m�I,:�|���"Ǐ�63���(�"��@TM�L�~�p�z�F�wb�IGD=�`�>�#�e"̙��R�W��P�H3#rP�A.��GXW�o�e��c#`BqNfc)�X��z����5�}1k��r����M�.f��L�A�>�R	�e��~�o &+�:n}e���/}p��<�A�y{�tj�z��h��9V����f�Y�R*F��}��2�3W�MS�A�
P�_�ʺny:�|6�E�����k�~W�4��P2pt��S)S�������j@ d��;�2Mʾ������$��%=��v�@�Ƥ���V�	�<�3�>"�H����Yk̙�@�EnR�\#˪Ғ�IR1�a�k)�^�����-������C�6�YJ��q���r=r]I�<���L�����Zxk�X����y{��9H��1��Lvx��_���o�38����_X3��zgRz��+��(pl(�T�Rp�Ϻ���������AK�U���=3_��{�7�a"�2�d}��e5y���l.Jz&ΘRB�U��'R���A��/��Z �@��m�$nL�B�#ʟ�s�\^����w�����,?�v,_�۵�[�D���L3���A�1j�c[��1�� �#?P�����z��i���������2xG�^$���-�y�=𹮻@cM3�f�l�i>�G�����y�����9G6���/A��i�N��󏛻[V���x
&cL��G7����\Z�9�Ύ9�'x����D�<�h�͉�)놵ɟR�dlJz~�,Xo��R���\J���� ���H�DF��p����!L���L61 Hq��8M�@f;Mx�����C�LfA-#ʘ��l ��6g�T8���nИd��M��"����`p��6?H�u���2���I���mϒ&=g&���Zp���G��TeQi-:�c���z^i�8�����>i �{i�y(��vJF���<l��(j
I�Y��~����}l_/�8=�E�'�g���o��^ڴw���X%�h����|<C�w�������5`��#Ɣ3��ٔǌ�9�ך[�֯��`o�Ү��&R�ѭ{	�f5�>6B�"�}�0]�&�{x����W��+���ȹ:/��x�)o�˲ ��`�		�klDL�ӯ�}�zO��(��$xV~j���`����/�%�c�j�>��t}'��>���)Wh�䲲�&앧x:0Az�M9z����o�6Ifev"c��v��T
���0�����{Vd��T�ZD�(��P[ܼ�"|�5��@޳��gEV�"�� HZ�p ã�ۑ��}���>�y�����J}�ج�
�Vi�U�Cy�,�S7�ձ��|�~�_�ɟG�q���y�]MGdJwۭ]Lĭ_�쵵Xo7�5�Y�����?{��������%���95P� ���Դ���[N�#E�������IB�w?�sJx�har�(�p���	�-��
Q�$�Na�ھM$�d��7�L��s������gd�=��f�����Qf��ܴ�_��Sc^�@h>i�5��Y&����-�8�/}��g��9d�0}ǘ|�Ã�����|�\"c:g�����G����́mΕ~2mFi�~Ed?�g3���{�`�������3f�($0�7��湕]�(��D��5J�_�=Z���	���B���	H����fƇ�%���׋���z���r���r���)��,%m�w����L�ӈ8M��@�>b]W�˟�����z��>V�?U�8D�ll�r�������Z�uD,�E�>)�MVcB.t�'�1��@���Z�<hrnv���	my�2ʅ�ZH{fr�>��j���g�.ob�c3���{�3m��?��?+��BM\d�aͤ�cҵ�����=���kG��>������nL7,|�S�x��2�oDm�t�����[��}YE�����ф�"f �oTz�i��mW{��}D^��kmϒ���:��+2��YiYۤˑfw�MnR���K@ʯ9ғڸ�v��Q.A�nn��#�SZ���y��ȸ�[%#�pW��ݤ�����ǂ�w������A0��GrO����
RA��z���P����Rr��r���� !������,�!b��X>�����O��������vy�e��:H�m;�dEO<g�+>�����',�	S�k��v9� I����K�;�����'	��'�V���U�}��z���gє�eJ�0�&�F��oˇ��N���S�̂1bf�I�8O\�}o^����sg��j�|.<�3	'�U6P�`̿7ݧ��Җ�k9ք�7J�<+�G������t*2o�1��\}V�X�(K���\�t�ːzud^?[Z �N��鋐r�R���'}�G�z������*�>秼���^=g�]ޢ8QL�&�X�)'%��:�pJfuR'++	�8{ϑ�&/�H@�|$蝄��������|��I��1&E�9�Q*���>%��X@��5&�/2���r���0#M��l釸p�>����e�^�+d�^��z�g�2��Li����u����;��̞��Ԅ��E��(Q��dIX-��0� 0T�ie���K̄�%n? ��u������l��5ykҶ���p���n�7�R4�`.���Jom8kݨ �:�d�����S�`˗�ᇀR�N!�x!�ibHU��uu��ȷ��u�y#ȴ	4��(��$��%s&�$��,�����G�\e��G�~��r��rE)���i0H���u6K��Or��,��$�m���%l���LSj��4վ���|���������z�ߎ9�BFa�%�x�����H��[���٪Vtp�����Q@"�z��v�N�G��I�t�����-_�~<��d4���������'MwZk�U�� ���K*�}��x%	b�yB!����tK�\x���W�sɗ3�!ns�����9B�%�Ȳ�c0�#�ܯ�����C~��2D�rw�B�f��|�z�c�kΕ��B�@� 3���ϟ?�:�����?��By-n��ϑ����㸙�Hш|���^�v��#l����j
�c^�٠Q����i?�#&�V{����Y�}�x�9s�%o�@!�!Y�eP�}g,�Z��V=p.�����S*�k�)�t �/�_� �?��q��H����@��=��~Wim�	X�63 k��f���c�eK���o�i�\�R���F�'!��>�ܲ�87ۚ��T��xI؝_&�����G��Ǻ��y�{�$W�r/���#��4V�Ȉ1�O���ǀXJU��ϗ�2�����K���ݦAF?cɔ7����v�,muDr�����}r ��s��V��_O���vc�Hz����%�-M���g1�<���S�d��}�$�rr��w�3�Z��h��L��n�,�+��+}��(�G����Hȕ��s����>+Z��qn)����=*G7i�n7�0��-#+YO*=�S���5N`����a�gh��]p�L��fL��_�.2LTy2C,�[?�e�s�������~�_=��k2�#G�p���?C��c	�_!�.�)��d���a�1�h*�Hp1��y��w,?~6���[L���7AL�6Hi��w7��$�|�]�M �����������aޕGP.��Z�'���PL!��H'zോV�[z��Ͷ��vF���. ���H{-�|���dq�l�����}jUW�5��������jf���H`�g(��ѣH��A��h[�.A����7N\/��s����1)�<\�K�=��:�˩��~�>$а����q�Vz���'ӥ*3��XB�a���w�1�%H'3�T�Q�#�<��D(�Q�����1��<Mʳ�p��ЇMNT�v��r�F��rZ�k�� ��5zng�ٖ��U�L3)S�a ���켈-����!ݏ����gd���J�ɟ+��~�O��������2'����N)�M�W���S*�p)���~ZI���ܱ��	�gb��9#��FR/�T�>�L����)�W�k����+�����n��̦[\���η�+~~�i�>\Ԍ)/����Fx���/01��d��.�F&3����ݘ��jK�ͼ|)�<F�??��k��1J������)/�����I/��r��yl������v��_p�[�w�%�땕k%T&Y�DN��S�i�u������-w��F\ھ�c����i#0��Ŕm��pH�X���;>>�@�1��]����%�vz&߹W�H����>�/�}j?�=�ӒΏ@��N��v��e�}��,BX�~�ޣ������6W�ŵ
hB��%����*����3������p)����K3��'Y��v������-�r�����{^�Q��6��m��S	y_獭Țd7_Fdy��3��BO4�cLdU��KYnR>�|R��]a�
�#�����``B��~�z���Q����ů_�`��r�V���cu��xDc����mX�/�e5�G�˟�i�Y�Z��d�}���&�^�1)k>���_�3���.=�&L���4�L�;j�E֗�3Qy�U�4�'
l&�G����wF8+�Zf�m}l
u�^5� ��޸:ۼ6����q��.�V����L�?C�:ۇ$<W�Q���[��c��WȱKc H�N�L	�(��G�y��4)ctb�KAm3�� �٭#�Q:��Ěb-H������iI����1R������ͥj�ܦd��X���Z:�At�ެ� �5�h�����|��d�:������6�[rQZ �ܝ?UmO	BB�0Z�xC(��\<���r��dp��46҈I�i22��ĵ>�L�ѧ$�2��L%��]bK8���Oy|K�9y��1+4������Y_P� ��.�V���������C��[���o��ln����ч�f���s\6�pDb���Ss}Dc~I�lQ�L �N�*��WJ��7�xq-Y�v��CaAs%<�q�,��`��-[�t��9�e~W  ����뚂�c"G���v�<�5�|.}���a41Ƭ����uY ࿎1|��,���S=��F! ������d`��H��F�<T�3�,��Bf��|�n��q��Gd�5m�~׏j2-�YB	�T	���SM��z�$�9�Zi�J��<�d?�g���I���٢��k������i����:��{2?-9�4Ƙ����G�z�X�c�H��� ���6k�.rIx�w][~v�ow[�9�n��޽����F���#u���˼���P�J��)7�4ˍO찋3̣��[L�S��ys�c J�(�'K>�dJ.�M��?��5��D,��h�_`���ρA�@
�!Jr�(_柅�ԁE�Й����B�˔��B��kǪ&c�`����8�Źj�3ƔI�w��������؄���|�e�H�?>� @@�����$�\Q��ݶ��t9��h������q���fRl���Ɗj&�Ou��r�@_3���j��`�qҞQ�o.�������c�q�A-�G@�(�A~���V����/^�E�cR�|0��<�X?(�A���|.�ϖ�sVZ _3��5ɭs[������f�ևZ�qͅC�=��Ӿ� W�����,.-��g��f�H���-�����qM���ec/c��N�r�2��6%��w�?��#�����Q3�I����ʥ�O�.K�1(( ���M@������~�������� ^�hҗ���;*n���2Ú��|�1�����W�L_���$/̪s��FWc�Z�I���9�X����YƧ����F��$ƈ�9�1+�J�W�Y��q@�&��/r1�u�/���k�`�m.>��
��jyԊ��mY��|��~i��ϺN1e3מ�9�VF����Ŗc��C� �P�u��s�>��[����]&b����FttJ��L���ͬp�kf�K}2 �5�����r_.,n��L���*y�O��%���m6Q�1f������L��#b�>`Ƈ��!|�92���/���8>!晶jR5���l ��d�+��%��M�C��K����]��wv1k1|��G��IR�?�X���)uXތ�ܞE7L>����q�yeb��b[�`A7��b�~=[��x��E$���O��L����>k~�\C�St���1[� 8<�����1��	0:kM����x��1ZGB�hҥ�	 %0g�Y�R�Q犵�%--.Υz�κ������Pјhs%��!oMad3+�r�x��H��`n4����\_7{]\.,���R�6�{�HT��M�4!MޚL%�X�r�
/3Bw&b2�-�v,���BI����^3i�M�y�:�mLJ����J�O�.&�n.-s�f��7U��>SzI��節��O��������\.�����rɟ��:�R��H��̋gXCw�9:~U��3�x�4�"���~c3�}�m�0��U̝]p��j�Ul�Hw��JP��!bY\�]���U���+Ε~Ƹw�
�Z��d��o�GX�qIX}*u�,9H��Zz�v�w�3����l|���^&֔��ǘT&���X��{���]�m �N�_ �TF��`���X�c��"��}Hf�l�NM1
?� 8�����-l����b���9\܂uX�8���\��|||J}]��aY,텷�'a?9[�J�Mw$}Xb�)mW�A�6y\j�I���mo�K� �G�ӂ��F����aƤ����� &����v8�WK�|�����V6���{�,g��T���}x���6����S�o+?���v�u�;�)�|�e���H�s���侞1���F���(I;����z�}k����o�����(������
5�t�,ki���$G��^�nKU���&�����f3���z�T% �)
��`e�{v����J�]oK_c�ݯ���_q���)�$ �F�D�Ȗ�Of�@�0�e�I[�������c,��\.W\.)�[��������z�1���?w��+�m ��A���˰���%��&}�����L����j+��\�IIIP�,���߶(�c�Nk2Y7�T��@J��6;�L[�SH Pw���d��Ӥzލ�Wʀ�~�]E��ד��(���?^��	SC���1��t����Hb��k��v��S����u�p���s�~�u-��b�xB,�ǣsv���K�wtR��\ȼI��#_K�ƍ )�)-�fy�;�ضNqK�F5�*��_!e�5��H0HE^�ƤXU��a��ۯ��>[\�5f;�{8C�2�4M�7^،�������B/��kr�?��|��bY��K갮+(ɪ1�c$��h�;�Yx\f���v7�.��C�.�K'q�?�ҿ�������"�����<j|����Y]����着�s�Q&R^����3'�﷕t��~f �]B�#�-�3��Z������~�W�㖵�w�ϙB��Հcfj�S2�g#U�kYD�
X�q ?��)_�����Ue�~��B/���e#�,%7�ķ�U'x|���>�L�J2vC%�"��~��ܐ:ʿ�_����(#ԟ�^�r�4k����"��'<��]7Ia�,iQ����7)a�hxڥݹ	1�E���HV�RHE�ݙ�{�)o�+���rs}애��͜��2K?��3	�]~�W/�g\����N0�l.*Zbg��#�J2G��Ӻ�*���}��q~n�Y(?7�L�c+�8���Z�SY;s�� \Wr_R�9�;Rʽ����g�l�%Ҳ5S�X3��-z`�6?���Z�ݵ��l�Ǯ�K���I$ �w�ß>~�/e���DDR��.pv��w�`a�����4�����c	"��I��)Ӿ �JJ�6q�0��v���.�K�)�)�M���j۪w>���Y��-�"�\3_g�3��zJ��%b���;3 �
���-��mQ�}����������E�yPX3�u������+�2�kj�I���"=z�Z��m\����Y�`d�.[U�����ޙ>�B����ۡ|r��=�tݶ�?����1�nMT�H_G�!+��s��g)��(�G.�=����G:���P�1p���~�t<O!��'}�9 �,uK�,,��;���
�?T\�sٸR<�F>q� \.�����1F|||��/ �۽�sɤ�1[nn���$�'C�O��b���>�Ζ�1�&�H��M���/��T $O�^��lϞ+`!��7�|���Z�|����cY\w����d׬1�����l*��w:�*�lH?F��:�X�lL�E�wZ}��="_�>��=˸�c%�8*�SO�=��[�G��1���Z�`M������)| �f�)=R���8p�1����{K)k<B�X(=�1���mr�*��gX�G�imzg6�4����u�}�b\y�smW���R��-��߻�dL�<��t[G�M���=�k7n̷�b��j���i�uB�l��6	�r������-.�\��'���L�쓹��\�;
��p� ��bkn'��D��]��q�\��C���0)XbM���`��3e瓩D������B�1����R���\�A*������w8:_�ó��Sb�m��r8�m��J�l����\%D��\k�c>��5�/z�:�e�����\�v}.U�\�,�!DP��W̱#r�?=}<JIC�яGdg�qc6R�8I�{:�%�氟�������՘b2�sq9	���w�,>??q�߫
����ȅ ���/����E&Ǉ�%ŏ\>~������f)��)oMƎwşy�(�0q�%��@'��gYZ�H�`�����{��ɤTi��R h)�F�H[dZ�Ιˍ�K!�� �E���י�6p��^�&1<=�DρO��u�f����Q�Z��':f�t���_�Mi��1-�Lq�;���L�Ă2Y�R�z���p�ɥ��s仝���d�Օ��\���҇{�y�@���{�}��p��n;?�Y�mȏ����`]�󬼢�#����eާ��r,׻�L�1ޭt$w'�ɜ-�zۇ2�S�����;�e)c]�����݂m�цѴ�ҷ��3ɇ���쾗6�˲����e�g��9ԩ��@�spK�zϻ�R�)}o`K�:of�m�9�'}�M�t��#�V��n>EA�X�ˏ,���
(sH�)�PbJ`���U��\!����&$�cÜ�J�O q����Uψwޝ�W<Ԏs�� ���#�FS`#��E���+����)�>��{�I(���x���Y��f-z|��:N�]�޼�n�I��w_�}g��Q9
B����\�@������m�Yi��Yϖ�7������s�){����ۦƫ��z�s~��Y-?�~L�����-���wU(�Ӟ�Hz�V.�ẍ�m��Ə����D��@!_g�ܖ��G���E
i�#R6���v�W�������Nw��)�"��)����p�0f������	��c�D�	',�9�/=�	� �5'�0��d|c��~Ci�;�f..s�w��?-������X�2�e��[���˸G�unL优&�g'�l��-��|�OS�k�>������6,eR�� ��l�����U�l������n�kl�A0�R�����qM���W���i�,b��}�-�>z~>to3`�����Z�U.x�mlͲ?R	�kh��1f�������=��⻼d����/̊{@��Z;��s����֗͒B:�����X�#:�ў���z��WJ�����gF��-W-͚C�Y���&��j�w�M~-�]Of�WK�&���������P��eYcJ�EA�˲`Y.�^��u��3�3b�UKt�&`y��Ǐ�p����_�W�����������+�#���,�F�)ߤ�u��	ɐn�Y��1��c���Y�L�4�����b-�?1F�~���S��H��TV��Z�Y[�m�y��'��g�Qw�̟'2�oS T�*���Z�|�`���g�RĥO!6��c�Kc[��Ƞ��	)8b7zl(���b��Y��vŋ�����n	�G`T�� }��ó��|k���2�RF �u��T>�~Ϝ�9�f�u�-P��x�>K)��ܖ"���!F �]���"}37s��wQe�6�ͪ����d�1G���;�Q�=�i�&&Ѩ��}��>��]�Ϊ�&Yeӿ�·,~��	�o�3����������o�W����_�ԋ�m ���5�ˊ�u��W��#x��7��d`r3�����q~�Lu��R��bC�w��f�J�	F����Vv}[2��d�	����)"��*����^(�LK�1X�-�x�%���s��nr�Υ�P�\biS`��<��l(G'F���ߑ�]V'� �WO�)F�	R3?R_%㻱�u	�Yߦ֦�f�V��� ._){�@Nі7;��Z�or]� �'ŵfW6o+O:��6o,�8~���f�����+~�	����6e �YY �+�ȑ���mʥ�8OaĭJ�9g����r*��/`v�I��t
�Lⴘ�G~�<�Z�
jۘ-]�o*����(��N�0�=��{Y��u���()�~�ɸ'��tK�������������o�5�>&s��߲X,�Ú���.�D,e$&�%f�\��Ŧo�~&����e��(�_���s~ ;�^�X�R&��v��m����,2Ėl=�)�e�[�u�M'e7�E��b�P��Z&�ټe�Dm���m��W�~���d��F�mQ�N(	�V���,KI������ͧ�;�ཕc-�X%A�걩��G�b)��t����B��^8�)GѿY��m���v�I�m�1�z6�a�T���IcM� ll��Eݎ*�p6[�3="�7��Ș�-0s�Xˣ��ߢ�:}������"���h��j��T,����@(�ALǒ�r�r��������Mc�9��!l�����������Z������{��/ru���:-��>>>c��'�������ׯ_�.��c]}���zX���\��m.�a�u	3]��\�������p�2(d��������]Zhm���`Vf� �қ}3���[PP@
Љ1b��|c��S����b^W�!֩�����/�1O
D1	�g6i���7��+��
@Ƕb�~e�5M�I�o�L$2f�#��l�����#�ߒ�VH+hI^Kn��XcFL.nb{q�1`]C�g���`\�{�o�\^��n~��G��������Y�e׺�!�=r�s���¬ʪ�-�m�`��Ux
x��=^:e�Q�h�(3�?g�2�%ѐ�45}J.���X�8s�\���.���34��c�P6��7u�Ճ��f�zhm;g��4gY�W~�"#���U��7W�l�MP˜rpF�kĘ>ӯ_%ҳ��<S���n�Jr�a�-�K�iIZ�c����=1���o�4�=�if5�n�v�y�}	�4ɎXO�;z��Z�`#�"F[�@Q&��)hV�I�o���V�����q��?�/��˿���U���z�[g�lʠc�=fV��w.>&����c�7��X <���5��}J�6�R|�:�>��u��R��-�4:�;��o�_��Hz�f)�r��~ĸ��;<��A\�_�:i�,c���=&f˻Hg�;4�Q�!���](cRcBh�����r��lRLˬH����{���*����#r�@���<�Nr��!���l���%][�>x��
�,ͥ������4�d
E�\b�J����O�cgD�^��dN�e`u�Œ����2��H�!~=��K�!�����L;�<���z��Ǫ&kZ�uk˞έ�,K��}��8�=�D;r�������owc��n���`�����,������̋�}���sO
[d��:$�� ��.
�ـИ��M,�<Ie����1�ck�)�wβ�*�{�����ń�}����1�������.�\i�W�vd��x�Z[� :�}��7I/uZ��l�b'���T�o�{�f�/�����1���L4�Za�i�ɺ3Ap�y����ǏFͳ�[)����i��w��T㟩���]R��5��Uuk���s�+j�����i珶��O��B ����ի���5��W��B���k]�ŭ�s�9���봶}w����	��hc�d��� W#s���$�I�H��&������0흔�tΙ�g��;�s��/!��3-my2�:���5C��/�1:��p�"�c-����~"ƈ������Ľ�Zޘ�ǀ���Jpv�`��	I&���w��L����a�|�p���kI�uŲ�
��/����O���?*��K�,��">R!}||`��CZ8c�����C[��	
[`;Z����<��1(��4x�:�����LZ����v[N���'��x�1Ouy�T�z��y��#pk��^��W���I^[$��?�<����|?r���xv�
��~e=3�K� Aب�g�;Ph��t��5m?h��:�i�XMndӶ�G�T�C�ܶ����_n ���+�׫m���;k�||4��pƏ1H "�����<�ϲ��O ���<����R�PyK��X��Kf�묣��>����cڹ���y��޻�9���O^�3B�g�w��yï?���Ͽ�ׯ?�0��dp"���vò�M�Y�c�v�lk�m;>??��cź����?�RI�<�.'����'��X�1�^�ޗ�\9��5���i��p"9 �%�-1Q&�Ax�*|���ER�\[P��E��%�Ѐ����98;������4�q���
��`�'��H�	W��c����Q2�#@�N���]�U��/�Z�������!#@�ujrM6!l7'�;si���e��j�mj�:�� r�Օ�I07|�/�=���nU�Mu�K��Tes}��6���v�Ѽ�yY��v����H��Ȧ�5 ����3ŵԾK���L&�s�Y�z�	�cY�[��%��\\��;�L�V�eY��� D�v[��z��W]��@�(L�;wz��c 7}�8�	����YB0� Z��mG3�x'HLI��z�w��8���M�zj��֫� ��L�U�<��yd0�RzjM�+cbұ+e�I�'�����5���<�$�.������&UOy�}XҜf����,p�R�����1[\f����0�_)@,ڙ�������t��j��3"Cf�j�"~4�z�	@�fZ_)&��\��� s���g�R�>��F�Y�|p�]�u���>&�Lk�ê��sI��DG�;����z�������~���wnK���f���s���Zj����|�0������L��	Lr�Kyxłu�z����r���%�XR�]q_%�Fw�}�r�'�+��F����,ȓ��g�~���2�
���1b͡vf6�3cI���@Sc%g7�WeVS�rT�;E۠i��o��IW�ԫB�d��H��qM������/���߱����-+�*�w�ථ��X�؃����>�r��9�x8�cYܲ��-��X ��`V�������O �4-\N<��D9��ΥPGٳ��Ź�	G璸�9u�c itD���\��0鱖�7g4"��B�a�����l2*�lb��
Ox^'�.�1vl��&r5����5>�Q�Ǩ��j���������W���^����ͪ�{bLJtP���}�}��ٍ�l}\i@�i�0c�E;A���W'k9�4##H �>���c�YL>�+y��~I|�6��T�8�z�JvPd��q���i�i	"M�Zc����'��yb۶�����nG�E �F����ҺS�-)�%@}' 16d������`���ܟO�ȋ�q2�sX�e]�W�$���<��n�� �4j�4�9���S��ЬPj)M��Z �y��J�Y���1��v��໯�+쥼��7�O�-�8����gw��f�� �;��.�`���3?}����'4��2fů���IV�h �W3S��;WD���6�\}��hA�?ԝ�3��� cQ=/�y���Lj�����y�̜u6�6 ��5���f������14!̨�����a �dg�� %ǟ����J��72����˶¯n]`���];h��Ce:�|��1-�.�d���'S���u
�]��A����ߣ*�3iv�m>�Y�G�Q�b���Lʳ��(���n�Ε�Gm���{H5����2ytnZhg�T�@�Y�ث"7g��q�U��d����է�U�^��A����<_��]x�	�V;ڳX���l�b,!�?�׆+��߽����3�B�.:KV��"�dz�h���E,��8�̑���8&P�<����q]������<j9ٜpIY��-����5�U~y�\�E\,��_�����@0IUް�Y7΂����&aT�	@yYz<��M�N�W�^���I���>�H�)8����be��ngB��,�kU2&�|���9M�WD���IM����_�~aYC�p�t����E��W��v�X���h2L������C�AS�xx�{8!�+&�y@��R����k�q��ȍX�ˑ4b���
@<F�N���Ʀ�l���}��\�#h��+7ٴ�*�#Y�u�s��S��#�ۊ&���f706�9��U�D�¨گ��jB��8�2�D
TD$f�d�|<�����>��Y7h�{��T|��3L��1��N�۹p�>�����?����>`d(�s�/o�`��yH��j)��a"9y#�t>�rFP��q�z�c�"3�wz|�+�#g1f�"��s�ғ2
�t�`j��Co�Wg��u������L��g���_:7��E��̾N�1+����:z��/4�^=�#�������B���!�׀����-�&:`��X�dk�:��N�,?�=o7֜�<c,τT½�>g�@�93�m+g�+�-0��^����񭙙�`����?k�.m!��4˖B'��6FX��u&&Jb���|GL
��M�#�ll7!���ܣ	�6 ��`C"Đ��k*#����\�sES�6�� ��ϩ���`�H�@�bE��'}�OH�
�c��q��� C���N�:�"p���N�3��W<�9Sh���|��&��c0�k�0|P_�'�W�h!��V���T�S�����,�� ]�	~��R�h�xt^�j�+����|5c���jϥ�����(Ƿ�)�ʨ}=��*o'�u���<3+�2�Uw��Ձ�RI&⁎{�2�ҌH:iJ5�lǁ�P�}�#ߗ�k��2h����������lN�o���0���x��,;�+��ʼ0�d�	4/�G� @����˹���$�;1ф���,����$�\S9�ԋ�P,�S��r"�ry�]�����#6���'�3|Z�߯R���]�\!'�Y�V2N<p?�����g�zv�?�|��/��V�֞�z��gy��F),+�Q�JM�+��p(�!д�4 ��|õ.�q�}6�%�������<�̅����+�c�͈�a�a����w(���4Y��>������ �D�Yd�zk�S��y��>`k\a	p���K>��%�f�}	p&�(���f�6��RX��م����L���̇�[�j����Q� ��삃�1ՙ��(�S�W�f�@��Q��>?@�j����-��2U"gW�8���v�g,��Ŷǲ=#g׏� W��H5���}�]_a2A��9r�9�f�@{��	��H�b/����*۬�)l���Qn��3&�u�cc�Y㙧FϪ�O}qv�>F0Í�,?rt����Zƽ��hg(m�.�]�~l��)��s�Ҏ�Le��'��;B)ޓ��  ��M�-�ƌ?9ĺ����pF�ZV�^�����7�"FDgS�hk�@�I���c�g3$U��[�U;�;����Ӭ�U愕����A�hg�p��	Zr4�2���,�0OIRr�v��π!PY>�eqg Vk/���o�(!Td�#P�S!���<F1%�ǯ��?+=6M.$�5�-�1svﭗj������yD:�W���sz�yr.�6 {��A���l�|���=*�׭=GM$+�Ar���φΕ�km��#F)��5F�TN�fw�4�5�&P��uy=e
}׽��>r$K���Y��i��!r�^�i��o<�m��7!$pĎ�9g]W����V3HW��/�3,K�խ�O���Z
�eصiN�>�a@��C�5"`�����{s���&�l@�����;�"��M 4��_P��#����&�WI���u�߹����14��e-��9���U��6�{���Q�^�����6^�w��T�H6J�	���]�.t̖=S�c���B�̀���c�\��u,����^��=Z���{��d_R������xv�ό�d�g��m#�-���6Ʊ�9��pV��O������2+G�Ɣ��Qu�>W2���*`�N,�Zkm����噩�1ι�t'�3@:"y����!nw�|�F΄?4ىHޯ޶�6k]���@�5�y-���:����#�lA�����:�	Z��F �L�\�:��w��P:"�q�q��+̥�͡����/�g��U��|$/�L�_!�A�3���
6)�|��Q�+"�9�#��?ϰ�W���}��/#��F�����A�w��`��ؤ(ć�+up��z��k8���aP�ڔ絑�g>|�I �\�̋�N��yy2�*i����r��45�C�<�5�_-��5r�Bծ��҃�P�gJ�Ep��Iӓ	�Ą<_�Mwb��|y�Ӥ�N��H���Z�_'o�lYM�`�Ή�;��2&g�
2�Q��3:��:�s�c�O�j@�X���i
���3�1��A�a���;�,Z�>^N	(�0���d�����%%�k&�g�.I�5k���̵`��r���2>�T�rf�g�ʟ?�s�.���me�$�p���\s�yd��UO5�}���5�OΎ�q@��=��^{$�8��G������,X=�=��hHr�;�R��2D���F��#mx�	�E�_��ϲ�W��r�Z7�ю˿S�A�ҶRW�k����F�(L)�������&��sS+��Q��?��T��V��6�Ε�a!,.�3��έ{�yC0� ��! ,�4�o��t�h�=�%od2#*�4��THS�5Mgk��%��l�A�0�z���?��Ē�`�� �E�[u�߱l��u�Y8k�r���hi�� �Tr���-��z�3��+ei�tn�>�yp@l��Hc�5�9$B
S�QrEo>�̩H�Ŕ�Z����Y0;cK�Ҥ} 3J߲��؇ �'���S���v��1���p�^}@��[��9xH�y���b	�����c�"4s�r�ꕩ�_+w���=��R7��P����&��qX'S�^��yQ�nt}/>fsl0��ĬԢmpo9'i���%Q����&I�u�͎���I:z���vr�5���X������'��_N����'��}��V,nE��X�M 6
�����%iV���m����2E�1���F�0��������Dd�9�:=p:�w�|~�#�t^���L ����j��J=�,������&,�Tp)[vCuǔ�n��s�GuG�4%�[�F��܋�(�v2m;��1��*q�o&\�#�@^Om�w�Zh9����v)�3����
G�ar�9)�إ]ٯj ��0�����Pfz��,XK���Pk�T�JV�Q�@�`���k�o�h�{<�$�@���3����P:D����{�A.�,�:�cO�0���4�6�g`�����ɼ_q�rno3 ��$ ~��x?�=v�1��1�3	�����J!�x��$���{�Jؿ�1�� ��ؚB��x#8P7Ʊgr
KFT���띵��ӌo���.Gz���Xo�u��s
�,����2(e�8���S#����Cr����� �*�\��;�W��W�H�Ϸ︠�Ȳ�.��c�����I���%l�surU�[.�
��	�}����[4����;.�Anf�^{���/�IM*^�l�&���ɳ�XSv�Wm�H�)��v_t|�A��Y&m$g���+��(h?�y���(�һ�lD�-1����9zN��\l9�Ӟ��t�ػW�w梕���R2�Sp{pV�u}C�C[�������"I��~Ǯ�<D]S���C��!��~߇�hM�ғ���ٗr�k��/����z��g8
K�Ʋ2֧v`3��S��W���"`l��і4M@���NP�j˲���s�E�\�ǽ�h7Sw����[O����l��PΪ��y/	����(���k�KzR���ْ���2��=v(d5��v>��eTR��R���n�T깐bsF�<�w����*o�z�ͨL�T�#),�R���z������賆M{]���<�}9/�Ug�U= J���~O�8�7e��
�k2���ikXƴ�]y��h�yx�����Y�WH��[�.jC�)`�#�8��?�'g
S�9i�(?f�Y.��d��z��BN]T2�Hi&�y�wy�a�J,̘�ڌ `�ΙK���P��T�3�$ �y�?�D�Gv Ĉm�q��X������v�j?
`qn��oX���3�9/��1�.�t��,Ù�����g��mc��cʵu�mz���v���Sd�p`4�|�N��弝1���^ ��o�3}b�Mjg�Ļ�2+u�h�T��3��_s>)��_W&��k���z[!���8�R��tllf������hu��"Y�YF���؎�n�K������k�2��h�\�h��π�����cp���3 cM��ؾ��K����*	n&d]����ﱕ�#���<�k^!Guw���W150�	Ʉ�g �-��-6��!ɫ]�����!b_��;�@zv.$2M���1�?1�U9�ڿ�-���k���L�-����>�'���	E�l���V�LW�pF T�H�ojNs��� �֮���>�2��M�'��������}��lq;[P��r��l5�	^���ZH�z��e��,0�^vJ��j���Ҳ��a����M�
s��m�Y! Mx1��ń`�F@tf�#��B\U��(��y[�s�HF�͵�!PM
�ڽw�@	6F2~g`�hF�R~-H X�ڑ����fv=�Y��~ǲ,�|�y�b4��ς���+�n�4ϒF<+=����_��9��eLfm�\���?��FX�9P򾭭�>{xϘ�͹&���2��o��K����]�7��3�#��ɐ��L ��"�Z��d�Ü�	vz����a�}�X�=L�%>�����Q]VO� �{|u��+`�2
5D���9gL��+5"�xّ�<������j�b�_�]:��C����{��10#RH�' ��ʊ{��r�1��
�J���M�ƒ �~f!�X/@�3��-#�O�w{��v_y��\--���1cG�ߕ���'����e[G��O�6/���5�71�&M��]��w�6��h�d
����EK;y�Ɍ���+8cI�_1I���W�9g����Z�\�7�T�BI3@E���5kN/gωU�Sġ�(D��X;�J�2����cL,Ⱦ���~��{6�����BnD1���V�H=�M8s&�Pc- <����)�jg8�� ,fDN�dK�S�{���$<D��j��Ww�2���R�BǆE�����5�H�6�8�c��*@����}����d8��~����r��w_�;���d_�7�2fU�tϥ}�:>��Zr��P�=�؀ɱ2 �O�0�vU2u2x>b,N:tlY���:�g������$��Q.�@*0��ܖ��aӒ��|i��ۖԋ�̉Z[�v���\5��[ʳ`��'�L5W�+�F|uL�4Bkݾ��I��w�)���nh�9��������77&%9ig�l�f������=0��������- 3ĸ����������'�������_����/��ض��43D�*rPG *$�N�=���@%�S]������F�~�v �2_VV��`:F��F4�&rG�u\�a{��c���� ��Z&
���fa	�f;X����Մ�63���)[׵8x�]- v�B5Q��IZ�-������Q�3�s�B(�W�"��hҽ�F�Q{.�w�(\�>�P8<�qp?~����u ����l<Dߴw��g��"��<Cx9���g���x��2-�����mT�y̘�ӫ�3�lS?��x�����3�����;��?/kB��>�"��3�7ur��-�w�����DN�	0���^,M���6��?d�(@������Q��T�l�ֲm�=����$�cAeG��~�վ�"p0�����#�mG�v�`���yl���|D�&�ꜚ��@Aة�ha����	������aYnǍa��4l�6:��-�6u�}�p�&���/������?���_�ޱm�m϶����!� 	u��������]�,��>�;�`6%�;��;���<�h!�<��n�@����������)Gt��8�5!e�il�$D9��dV�^[�)���9�K;=�������NH Dm  6��h��gҸ�m>�1�⾊��:9�ņ�o|��>����^h,�&~�,�ƴ�.����jCy���z��c0B���F��l�Q�A,4�|c�78�v47h ]
%P0�\����_!rs�O�k����ןm�z����#�ū���|���b��?�O���^��ʣ�#]{�5pȠ䐊�%L���3��<��9��-0!"|�۶{�6�XC Ч��{@fLv�>�����mKw�m��6�#�b�iк�� �.޺��B�F�f��ܲ��_)�E�����&��@̏
/�Z�G�c:)��fOe��� 8�^@v�z�l�\�ʽ��.�/�M��y��'q��fd/��S��0Vx���z ���D��Y�Ψ�볬�(fk�NU��/`f�4����=����=�&ׄ�޴���:���|��0h@��i <��{��SonM^a�{o����6�W˘�����!�q1�NkM	d��98%��I�!�w���l��e�~���QOVB�?�c�	OH��m���]3�%���}��dF �����'�����!���m4w_rt1���g�{e 8�Q�տ�w��6ͻ|D�s�R�uF�^%��w���A����w���"�m�x��pE����/x��	)�ة\����w�<3D９E>���E��TY�w�������M(b����J
�C[2�,U����'؉���؍�@�\8:���l��F�XS�_eYx�`6,����m�WK�^7��]��Xc�k�y���!��(=!t�@1#����+"�f/]�Y���?*�~<w�5ǜg@0�r<j�Q�>ې>c�1jo�e�G��qY෽�'>�^�~���1�F�,m�خ��W����O^���a�v�ۆ}���p��x�7/�&*��?��`�]|�୨/"���>��1xU'�4��u��h�I�vU =˥��Y��ӘcV�փQ�j��9��=̙ -�b�/=+�G�Il� _�CQ�JY'?Μhzm��s�3t�/�Zr�։��r�ٍ���D�F<*M��2T�ֆ^��jt.�B�1�ƈ~ǎ�zG�����lLe[��H3��A�0b���G�/CSOS=�$m��䙸�]���t3i� +@Կ>�m�Ϥr���Ɓ/�Q�A�q�n�E.#a�{�v��s Nz���/tڙ59НE{��:�nsܶ-v��^+��&��	�l!�A۩ā��e�|cI��gV�̓,R�qp�pd��}�G����]���(�u�Ȉ����猼/Nf��"����,C��YA"}J�������,�i Ƃ1�I6���c��#�#ϡyF�!yo�ث�L�9N�z����������w�qh ��uZ���9M��ζ�Y�\���9 �6�6�u�"�y��D1��c�-���;m= 6�����
�=�����¥�ʛe\y ~@g�e��{dzF4�%# p�Yl�05�?x�X^֙Ͷ��<8�� ��y~�X?�do���5S���9�!��%�k�θ�+|�W�u�qfJ��%>9���g��������IW�\�gm,�]98���1��\��#��X
¾��Uw ���CƸ0���c*��٩C��	�X|�MfwG��� �\z��MDe=���.:�g���v��;�9�j[ǻ��J��q<eH$�m|2��r�8�1�c�C4�d�U�1}<��bBC2�f�L5���agF�8>kw�դ�(�>�3��Rx��Xg�0<�������e�y;�V����|��T�G�Vf�/��>�=�չ�1{�+�~>?$��+��g�#0���#5��,/<h�9��&�$ �'�;;W����v2?[�ɻ<�i%bkj#�؂r�,D�����O�̋�i%c��,���щ��g#M"0�~,V��ڣ��/[��1	��ᢩ ��3���l�J�lY���,d���P���/����2	l�͎�gj�u�hǩ�UgU�i�����-ڴ�Kol�ox©=Ze�j�<��d5g<����]�����=!F,���`CK�����=���-Z�4M��}ɸ�#��:�Y*̃�J�.�̢�I�3���c.r��E˪�H�	���yM|WBt��0����Y	'��Wx��n���u�C���I�$GO�g��� ����q�I��N�?�I�! 4Y|�f�B}M��-o�֎�I�2CH�e��CM Ę[i d0����s[gˮ�f�9��Rb��1w�@�+?���n0�Ѳ�J���P>N6����G��:��1���״���l7j׮+�~��XvW�Lކ�}U�a[睎�־�rl��;�8�}n�N�F� �ѷ��1��1<s�v�@�ؐ&A�#p �1F|#�C�k�m�x#���/�aC��Ш5�]lO���Ќp��)K���m	̩|������<�:�f�י ��E_ s.�cM�5��sa}Zcz	�J;�MO�j�%��� W��K[���0�s4e9Z� �ke{GN:W���p��+��3��6N3m�+�xDC�{e�ϏƵ��=v�4d����FJ�2���& 6b�X�7���T!�9��`ҏ�(ȳ:�}Ç���x��!3C�����+�fy�Mf��$��ր=�d�#��~��X�uISJ��'Z�wy:�	��}Ԯ���{�N��:���v|�5ƒM³lb;p�ݕ1�dL	՗X���~8p៟����M��+]���.�I�Q��&�.�8�m�R���B=!f3��\ή�Ƥ��ʌ�W�g
�ŭ$��Du,KE�䆋��9�"=jo�3�f��̀��Fepfw��m��{smv��*�zea���t����ΏH��Y��~�!�&�Ei�M���0���bfN� �#ܳ�<�����{oI�l]u� ��H4�eW�^'7�1�B� %x�=���&�����3��m)Qw��=\�����1�t�����Yga��1�%&�9F����׉<ߍW$7Ѻ
�N�H8�!�JN▩�p�*c��7�
0-f�+"�8�0�s��⋵aB�&�"�������y��x��� s�]n��Ui�H��&�1�ʦ�ӈd ,���Ѥ�6�}�	p���"���ٸ"� 	�AI�5��S~L�5��mLb��Y�(��U����ˡ~�:����{����m�l�ū��LR=��ůd�y��tfy�����F�ڃG9�*RC&/G���g�§wcxV�Ć����y��b��8��I�2�����s���@V!�L��<�Ho�T�S0��~'��-M�b���ΉLz�ܛU^��}�;���ytq!�7���\~����GD:qժ��ʗ��!�y)��j?���}+�ڢ��4c}͑F^?#2��hb��T��ғ�!)LR��.�ŀd6B��6���Zxkm��5��I�R+O��饭<[��YiTv��q���L40<��>�t�� ϴ�n�.�B�l�
�<г����|��&nj����p^��f�;2��8��φ%���3�g���<g��ks`O�m�kҬ^���Ek�y�C���e���ٵ1�X
���1��oe����E��i �e���Ǻ�)���X�0�U[̬:'Kڔ*�>����˲B>e���c̆�m<N�`���u)e�Z��왫ߕv)�<�v��O�|e��������B�8��Ҝ9Oc���tP�?s\D�D�;�ԝ�ZV����6� 񭜁�n���׵�Z�-��5�d4Ѯoԋ��_�*�Ec8�co�}��������geH�)�?������{�ۉM�zM��#��F�i��ֹ����	�k�5���93�¿
T>R.ߠ���jv�=���vds9��a��X���Z���!�qn߃�e�����U�|cܮA��}��1h�6�t�엽y���<�?��Y�/d�m9�z먪Y����ܽo[o!�N>x8��k ��ȸ�@�/-{�l⍁���.X��[\�>�IqsIc�^��L��7�{�Lc�~� k���uݰ�+V�/�u��!���Z�:EF�&��~ڑ����ɳ9lj�`��1c\��	MZ���"7�J�^�sG�ɿ'�7�g�L��Ӏ�$=ε�չ�L��n���+�4�O8�mfM���\G �6W��ە˙�W����3��s��@��%9X��C�p:=��\L���-������f�܂Mq=�{xY���&������0�ܜ��ؚ�����H��Q�,����i���r$�b�8�������$�b��hrmF���	m����W�W�����������h�y��h�f��y���5���7��h-�uC'S����޽x�s�� �������˺�`�V�e������i��5��r������N��|g"�����Y�!�99O)P�P�gMڬ>�
�OL<�e�F�����{�B&�gr�sy�Ʀ�sn�^b�H�;��O��4P�3iGV�'�s	*%c+A���<��;����3l� ��N��ӣuj�L�%p�#�&�-��t @�[yn��1����9�m�v}ڤff�|�ݜT�5���|Y����;��.��ǅ1����$��6x�h���t^���q�=T�W����Nj���k�u!g���S#d^%چ#��98���[�A�4���}�9)`RqP����!��7�d��a
�� r �f��A�2�Y�~�e�aU��I
m�&pi.ˤS�K�4��w�Q��@JPx
�ԀGi|>�� $0ʳpFD���Y�{�+ի�����{����1m����߳o��"�V�ʤ.UN��xf��b�W�tK��|-���l؞Q�Q���{~�1J�Q}���$���W��/-��)�"�\mE����S��PG S��z�A.U�=����e�F��T��t��rv�rU�Y�10����X7b��/��f�����qEZ:^>�'ǥ�nj��*�Q�h]$r�1iqK����n��2���1���ჲP�#ڸ$ƒJ��u2�=�Yl��C�9��#d�s�aꦾI��d.+�_rq�����-�;C�4���	(�<O����:簇�����l,�����J3yǀu�(���{�pY��#k=F[j��NڿH0+w��ݜ��K/YZ,|P3�z�>�6�ءL�L�j�cL��X����E�I�>h�J�Y�8:��&�E�QnOŁM)� �v��9�D��A�d9�\��e�(*��Z|�?��^��0ƨY�D�uy-��jGfe��I��4���3�e�#��דW��ƃe*fyMl����EJ����D��:bs*[�Tm��c��k����<����c���g:F�J��g�c�/3M�kW�N�Wg�}�x<ڈ��@j/1�=�6�:��06�g�&}s��s;v����dU�q,L0@���嶅nV��)�񶑼��ޛ��7����$	���ߋ���F�C��Ȧd���vKv�!`��a�$�E�4���`����l�l/��\���R�^�za�NS~>S�����j�7c�;T�>�Ʃ����H�/�h���ش3�ǫi���¨��&),�9���^�����y��MG�Y�W$ƣ�4�QN�<x�V�l�bcI6��y�ڲxͼ;�y��l���<���=v�U�q�ܧ�ą�m��$;�3��Z&͋ϫ���ڵ�G��V[��#�I�gM4G���$����!�믔䘜6����!������?��#L��k�;�9 ,bp��6���̀��@�A���g��aY�}O)�l�&�)"�h�\̅R�����(�Ř;�95�x��y��ky�i����^�"����Ak;s��̬��]��N~�y�<��K��Ef�>�cݝ��:��W}��.˓(���A�\d�ϫ�R��Ƚ�s�42I�Sm��:#�0fk���bFm�j�G��\�#������jY� �X�We�	h����ֶ�O�窉��\v�Y��5V��?}����d8�1�-��C;�Nl�N�l�8�Ҽ&�w�)G���m�B(�{�Ou9	C�.{dY�8�8��Ѩؒ~�Y�)%Uy.���X`b����P@�ӷ��"[��#:?�P��{2�	>��{�M�����'��4��N�hp��x�W�1+)��ya\}�v����m�P!��. ���u9�k��;���/$�)ck0^G%\O�k�`dj"ձ<D�a���1Ɏ���mzNN��>
b5������d�ɛ��g��3Or��{���m�����3���g������͖�d�|k$�M�Ȍ1��i��$��k��m�1�f۶-_{p����ml�m�#!=�}ے]��Ls$N�*��]^�K-lVAX��1]>f��jh#���iLQ�c]V��{����<���烢��j��(���.�h��=HkKB�#�#/�l�9���츌1�}|�n��f�0�F�m#��wH�6�����h�s����\�E�G��U�]�71�ϲX���l�x����w�,�g/؋���^[���#��)��V�<���H��n��x�)��-uJ�b�J�H�P	\j�2b�T��	�rַz��C�������Ӝ{f�.x�(�L���qqG���2�0[Z˒��=�f�	m�%8�2�mV�k{�@��+�kF�#~��D�#����>�ۆeqp%�r~>�g[K��!V"&Ĉ%;B��g��E�N!&'���Z?�,JeN�η�[m2��B��.P�Xz������N��F�M?� ������߱�=Ƿ�,>�w��/Em1����UW�����Gv�3Ҩ�Į�?��d�ۡ7u�VU~e��ʦ�M�9��yn�.Cƫ�jR�أ�t:�^�%���B���R�����y����Bv�@gāe��W�j���+R���N���]��l���m()鐦9�4Lq�Y�w�y��krU����$9����y�*�:�wgʏ2�h���yrn�i�f�6:gdv%�	�:�f�nt��Y�4�&��c�C!o��U���$�xut�$x����O��3�J������|��d���c�]K��G�k�t�';���%�� 1�)��X�K�zJ����Vq1�4��ő����W�̊Dm�@m�!����+oV=���9����Pr�'�:�=�b��Z�	�1#\�~�Gjy���r�x>� ��s/ߊ�\��5��v�-	1��x�"�E�K���Xoަ��v���VX��<G��"�U=7sЬI��
)�(�<���V[�%��#�<�&~h�k��g�u�6c��H��asV4kyL��d�7��˝B����U�L�°����7��2��XS;@�Y4駲���$�<��ɅdPi���afr� �Z�9,��, ���ܖ&7K��L�z���t�g�1��'<|����zl�Y]��[F�Q9cxϯ�9��n��x�JVMk��
�<�g����H��gm�YV^�s%���P��̦�C���#m�ﬗ˜�� �v�<�M���p�%�U�PB�ɶ�)�dߩ򘭋ͯ��9%='��Z�4���D�W9w�1X9I�5K�YPy�z�rif��߲ĀW��e�d���ZR��u����G4�r^�w��I���Lm80�_M0=+�S�#O�HJ�1ǯ"#���l�M9�P��x�8�����f#��6`5�$PgM,v���eY�-�]�T�S{4	A�`k�`yT�l[4u�TKk���j�R (��gl�<6�7]���寨�f�?g���{Q}J�=*�j��S������k�Id<L^�E��t���G,|�qٹR4��������J�3��$�S����4,�\\��t=��Ce��(8�������m���nO���T���׫����g�k�9��mL�<�^��i=�0��\����ׯ_X׵��<�	�[����\��m͢l?֢�n����Ʋ�?��)�|��@.���n�>h�������)�#R��u���_��;|�����Vũ��ް�k���aYL&�R���.�������pR�������p�o���0*�:C~P��T��?&��թ�:�/��-�D�Ӽ-7�ˊeY��5'�O?�{�"*�<H�S��쑌RKʁ#�`����.��c|�� ��J�l.��-���y0�H��W۟I��U{N�9���
�:��Y������_�ʅPL\}v�L��)\�h���O�]T�/b�fB,�j�||& <��x�Ş�b�A��^������U�e�w�Y���l�J�9�W�t<�ˊ��,��=�y,��v+,\��ňn���X��>�ʹ��8���뻄Ɖ[��β,p�!�5	�fub� ���+�κ �ʾ%�-F�H� �o������;�4MmPT�+3�DVE %�$� 'bD1��h�C��v�C�2Ǝ~��pyG��_c��+j��¨1���Wv��v����~��_��L�O�P�@�����@�G��Uu+���
0��ۋ[��pO�.�gm�|���͖d({m{��'A"��P�;�T�a�u9��2���Y�2�09��)Hɐ5��_\�:�Wߋ����Kt$|<њ�c.�s4�[2�QY����VI''��Dl�f�$Fԟ'�Mx	 �	�f�Fuy�>t����'��)�db�z��@T�hgS�l�l������c�bt�X[�dw�!:�(��8&�V�4/����>�,�{ei@����Q�����-�j�ٲ�I�O)Vg[���U]2����&r&����Y@xX��2lϰ���>.ݾ��	;xY���2�e���<�UOz��IA _m�����F����h�~\7��zh�5�;V�͙�G�J�%Wڧ�Ui�f�5y�%Y��:q��Z�|�m}��c]�&$_��Z���Й�*����ݧ�<>�}4!��*���('�F$�[#�rgj��Η��_����>u�A
.�Z�?�9D;/M>&�E���Ͽ#}cҧ#��Y���C0���,��"�M.O��c��� �k��|Ѯ���e	"�/CV�1>p55�vO#{�]}V����;�.:{�DMe����} �k`S;��ď�\��MP�Z�F��w�c_�������Č|@=e�֜V��e-y�����F��rv?��?�Xё�����m��w"��wM�(g�u�3G ��S"�?.t�~����w�e��L^���9�֖\Ρ�XͺJ[�ګ��{s�F��y~�������$�	o�I9��kZɦ�����@����݈?#����vYBHi�?>����������o[�|��ؘ����G��d�̓F� ��H�W�1s��?���m2	T��UB��'�ʓ����px��s&�ǈp2��ˊ�-�g�%�Bq�s�^;�`�Ŕ�8�����|��Bglg��ɧ7�\�ݾ�_u�,G:��3c��kz&��N���'�g%��?+Z��X{��}ic�1�+�����)� ]:�t�{0���zޟd���s�(�U��`[���7�jZ���f�ƽ8�p��4ǩ�C�N��6�ᶇ_!�pF2��z�U&S�UD�p���Zs��٤. .�֎�\I��>9�,�E�ےf	&��(Ƙ����;����"ϧ�;���O]Nh2��1���
6X�(q�J���eY��k���UK�y#~�M9�	��{EL��r�Iu0q5�Yڄ ������)F���e=0gm�Flb��c;�q��H�&z��3 �1�P�>��N� �}Yhl��}�^�YR4�h:�Q=��C&��G�-��6eُ�K͟��h�yP�d��[�'�5�=�x�QR��6jτG�Φ�$��g�Y���3����P;�旯]��5�{��*�����b#�@�����=��{�c���.���E1DF4ǹ���a2����;e��1�>~�+oa�T<��)0� �j��Y�6!��r�{�DD��I�}�۾a������??0�ֶ% p�^��c���=z9Q�NF^vtN�	��A�ɻ?A=:1qp�Ni��'��j!CdN�G������|�͏
IC�Ձ�G�j���̂��F�գ��\݄<�LQ'��Y; ��X�B�o�Q:�^{��Ng�������w�4)ƚ1�|Q�|(��#�ز�AF���`�k��D�h���>g�Imjߗ�G����3Y:���{��V��ڷ��F!��˼Ft��hs���p]�l�T��PP�u�������1fЈ�w����M��:�56�H0 Й6-�۞�#=���d����`��b-ܒR4��j/d$,M��L�Yd`\��`d�L�'���r**b&%�/�ԪR���=�/�8���+,�QM�m�;U9����v\UW����U���f���A����L�	"����iX*�fO�QK1�4�bd����X�+=YOէl!gR@͉�L/�h� �ԚbOi�v�+�_F��в�g�M5\�7�l�yӛMWG����;�s:���{�gg,�wB����u�C-8:�����#M�x�
X5;z�C�Qy�jI�����f��%����|g���^u��g�[�����r���>�������}�����W��	2k-nˊ�⟍�%��� gm��W�	�� ��G���7������Ox��<C�^����K�h�6��}�Ì1u6�cG$g��d�*���Q�5rw$cbg�3p�,�HR�����NB���M����y�[�X�H�¯W�r�@���"Z;G�?Z�C�����;�p����X��z�<�sO߯��X:Ϛ;�TMɠ�/|��V �&i�cbҏ�1?���u-�S��e��x��v�=3��6ಬ���Viï���<�^F�c�b�J$��=���M�����ߏ���)��=~��hG�bc����#����=��}������"(s�?�J)$�Ϟ��ƚZ2F�<bk�Y_�)�%~v��XWw�ָbs�MlM��d�ɖ���\*���	�a��s��JJ;KR����o�\s?��C�T�Vm���ms�6�_i�ܽ>�`<+�&<���p/��Ŏ����fWyV���g�����֖Q��m�^��6���=) �s������Z~�����3 S��U���<_�ՒT��f?��UE?�6m~$�� ?~V�H���?rJzt-!�Tj��Ȏ���lli�#҆���;�cE˲�'=E!Fu���䬽��h>^�IX�X�0�'~�s��؜/����s���
��7�q� Z�C���TO^\ �t�@�����3�>�e΀8� t��9�9;�h����ݒ�&�Q�MN�C�b_��}�<�Hjj��Lh?\ɳ��
� �����'@�[�-֏8�|E���F���B���S`�L��g�Qa���s���C+=�S~�y�w1y|> u/�1i��J$�a��y���5p��;���VrE�����kF��9R"g�ǂƂ�Z���V����,d=r�r:�����$<'̭�[��d��l�v�!���H6�г���`�Ǉ������-�s'��$�̰�D��Є�cK,f�Ǡ�\Z[�9 T�Q�c}>���jpM{�3�4����N��w�R��ULƠd���jDo��fh�T���?�*9�[�Ю�����齣}Q-��U�t61��f]�گ����!�j1�vv"��v\ʙw�3Yxg�M���T��g��Ս�u}p��{���9>āP�L�7㠣�W�}TF�
�&Ve{���i� ?^ݝ����������v-�j[{���Ȇٍ6��1��5���#*o�\�h�d}R#ƿ�|���ت:Ьu{I�X�HĈm;njK��XP��=s=ҴJ�iL�.�\3U�-_��5���(�s�i�Lֱ2��1&z�9��X�7����p�ƚ^F:3�Z`��]ܥ0�by�U�u��YK�fjӲTS͞���wb;�v���x�x���U���`�1C��>p�Ko�-l��%|��H�~L=_q2����2�6�|ϝ��1%%n�|�ny��^X�GU��<�ƞ�(�U��J�2���rў�>���:4��g�A��ӵ�����T�W��i�[_�T���x���o����������fQ�eb�ji튈���hi<�o.���)#`�L��,�s�ᴂo�7������όf�X��@�P&?\k`b����hdA� ���@� 0�G�+j���?9���D*��	��oó �����jm�l�OL�?G�Y�:g�������wȁ�왈�B�Je�� ���n�"H&��3�`]l۞�[?4�&3�
x!��4�;g%��ՙ#^��1'8!�ڡ�iE��Y��~f�ϛG��L���\-Y��h�M"�4[�U��W��5�\iO>c���k�\׵���bM���r�G%K��$0'����[����!oaD^��L/�#I,�1@��>��3��#�<�O s�;,�h-V�Z�s�i��:�L��I}X�fk�)�R�h*R�c��G��,g�{��=�T��1mA���$C�kcQ]vT�R�{y��`ӓ����sf�>[|Q��ߩ�n��,�����O�$���y~㡠 4���N��jt&�RiF8�Vr׋bTG�g�^ z��
:hH��޹W�זw9i��h�۩���u��ɤ	�KH�ck�kC����S��樳�>��9T{��s,[��ڊL�d�f��U����
e�P�s/�ބ���� &�&��y�� �j��M*��)�� Fχ	p�I��[@��Ia� �4XR8cV{�m�!�;L�p�)AL�ԟ �Z\�R^���Y��jsy|��>��Hӳ���UI�" �w�X�S�P�������=����!r�[����K�Ǐj+e,����f|��~F���=�g�{�Rv��9� ɉL�������'�D�fQD8-��>
%[��^�=�����5M���mҤ���Zm��;^��ޫ���|/�Y��H��MLmu���0�����K;�Y�P���WΛQ�j s�f>��B��m�M��<H��5ψ����ŏ�?��  �����ׯ_���ݫ<Ν�F���M�o7j�~��s�$t�7�Y.ρ�^� ��K���nXn7,��R �4V`L�X�L�?�� �����?�� BX��/3a��?19�$d�zJr�����"��;!L�QDX�lm�[��ѤW����m��t^6��ם�4���6;Y�@�b�s����	��qnwb�@ju��(}��n�ٰ}6�r�Z�K?Z9����& �"�*���vY��U�yR��b��q��m���h�BWr]����\���0_�	��oyǋ���_�,�Q�Տ_ɰivl�zf���wI�,�}�}��d��>*r���?"g��e2e=R�FN��?�k�l[�,K�H��̽j���(��}KD�y~�J�����7Ǻ���` �� r�%b��h�l��DcAwm��W�ȵ�M	�d���O�Oț��`"O���LƊ X#L���& k#2TE��\��r�23aXgӏu)oy��eElJ�Q1������\[�
��X����w�=��M��5����j���٢p��� 鳠�_n�A	♿���	�b��5[���6_)Ƥ�. %�>`e��~S��Q�fe����=�c$ �����:�R�J�a	�Sz��eR��W�+����l�O��V�u���b�suD��k������o�	e������&3@;���ߗ�a[v�9LM/]|���R�2cL��ɻ��2�-%��<@�5%ES��� �����8-
�)@IC����G�!Ҁ&�7;�4MN��K`v %-��t�1)SQ�i9>ڡR�2~����`a���#厄��~eٵo$��}K��\e�U��s�R���G&mcBI��c(���H&Qʌm$gDi������Ѧ􊍩�W�x�τ������E��+`�↎�u��Q�<DF��=;���Z��vl2{������y������[�vK������s��ͳ����}|���tΐj`��=
�I+�'�������=���=�h��1�:^���3;�J��x�iQE�;f��?�d���L����DM�?��Z,n!Е��L�%�GDkL^tw�;������Xc�[��c-��.�۶����O��X`VG��:����;g*%z�ڷʬE��Ui�Î/��Z�ib��&i�f׀^�<A/���w��Y�g����>ҳ�]��޹1O�d�����{�S�Ug!�a�}8:�H�w�Q��l%c����uuoe�x
��wug*����]VG@=.�z�����'�s�y�&�O�@�I�y���P1�=�U��!g�{��k1��ԟW��i��9T~͘�G,I�;��δ��d�m(���<�y_uM�2�4�A� �|�u��gW޻|/�O��eI����m߰��u]����0f�s�5�{���ö��}����;��;Ƥ�5/<&�d��gZI /!�|��?�E� ��b.Q�DcL�י4I��Ƶ⻬B�Z���.�D����n����	��h�zp�F�o� u�bdOC��l>��@���@�>*����`�l`?��|����@Nڄ=z�W�&+���yt�B�*��U=��<s9�w33vW������s�x�,�AH)$OC�\x&��j��ϖ�Oe��x����r �O>��&��M��֩Ո����ZZ��o����d]�r�	���v�9?9	�w2��Ծ}�J��Z����1�˲4�r��f�e�Й��Njw���1ѯ;`�{I�����e���C�b�L�&� ��� F�<��0!�f�^��D]��Y��N�xN�i$5^Z�W8k��|��
�y�
�fw�V�t\���d�7�+ږ�NR|�Jer�x�4��sfR�[�Z;j�W�ɵ�e{
K��ܞ��W��vc�;��E8�c[w�u&�w Y_%��f9��cB>"lw&��ԁ=饂Tϝ:���I{<ɍM����Ŀ/�3�H`�{�ኴs�c"����4�u>�1���(s�+7Q$r��hr*��sm��9�6F	Ɔ��j�Y2�X��y��#W���%jL7A��}҄䍂s.�@���ڽ��$���n{����K|��/�$����w9��A�Nd���|���e���7��`*�r��Ҟ2�� �k��s�0#L]-U�K����Y��8�`��|}0���2�r��u]K�%	R�D������M���Vz��W�;j�l�����j.n�xؔ�R��վ�l��BF�cΘ\R���B�L������"m��m������gFs�W�vo��Ѭ�m��k����Y��H֌�Nzs!�G��5@G�{m�>@H�ZƵ}~�FP�)]5 ��Ie��ہ�m��g%�\�\�4���j"6�_��GbM�� P1D�C��f���i�O���-�6�rb/�G82X~�Ӳ^��N�1�IUF���^�AO�cj¦	����x�����|����n��ڨD�ۉ1!$���&
m�xe��O�=e��;j��e8�v2�]^�M�x�����|@�Ύ����sՆdX�}���r�ۻv�&�{��Yk�>�vm|1=2�31�=��LF`X�:!�V�6c�&������+v�)�Cٵ�MܡMY���<�~n�ڜ߱��6�����s2w<�?��U�4�ÿ������g�Yۥ;F�0�Ϗ�6_��5ђ5���|Κv�=�k9X�㷏��U�^��h��Fmi�zs1x�H�s�N^'y�(@uT���R{�Z�kѰ����z@�|�Q�1���5p�Þs�S��4��7���h�)�]�!� �8�w�{�m5��Mt�[�-�= 3�35ye@��_f�V��ѤRHLc* �4� @ ����;�}Ƕop�k�z F,n��`Yה!#�n0���$g��H�ޡC�l��t�=5mk���1T��%�[=�m3Ip[���0�@98M������O����g�����l�8������[0*�<2�����}����cv�6}|7�$󱓚q�|��嘓��׵jn�1x�>ٮ��)��Z�ư���f������9�G�~��q��[;�q�R.�kG)�0�`����%PE>�3����B���QX d2��sd��I�Ƒp�H��C�-�H���&���u�K�ɡ��P��"9�dGhg�1s��=!����!��7(9����mJ�5�DMr��6g�/Z�Av��Pr{ҏ��x��#9��<�%�x�g�=�Y���y!x��G�3�����/���1>��␓���0�N��ֺ#��Q@�|�����,4h%���u�u�>��:�+��U��i���d8�|��`���J�6�I��3~���Я
g*yu�9g��J���R^���9t��7g�n����~�8�Զ_믜��cMcy�#���h��Q���v̴��B�}9�a<���C~��t~{�L$��v�J�Եg�,�7\h�N顯�d򺈈�,@�Ԑe��_���!o���>`π��d�,���K�ͦu�g�-F���\����t�C͕`�|�eI/�&&���ڸ�$����S�c�������umʗ���>���c&IU�'���з6�PX�jc9Z<88��������\���'�4)ml�9���^�g��3�C^׶o"[M�����-g��U3��W�/ύ�<2��+3�\�u7P�G�W�5�ÃU7�3��:�16Q��(j�+!�f���[��@�b�`J�����l� �cM��<h��y�|�w�/� r.�D��{�i�*ia��w t:}Kf�k��޹�����r9�o��|*4�?+����(���D�U�?�(��{�M��ݧ�X�ߓ{~��I���%���ʒ �
�E4�L�VL�E�lL�unkjH�!�]��֌>�����T�sX��۾#� �Ԡ��`�F���;t�}O�zʊ��� ��^�@��=tr`h�}���p;���&4/���L�}�����r<[44[������uk�֎��+��G��m_�18�S/�3��ɟQo�t���L����	
 mõ����Ҧ���W6Z�಺�bh�!�4�^�{̣Yg�K�Z�U�OF�9%͹G�xfn�����c�/9� BG���{������̯*��"�i��B�ϯv�5�78f����z�Ck����v�!��_��j������qo�նmX��@��7��=�����;vo���C��c@��9�������`���=��yP�
7��'���-�l���jb���|F$���2Mƹ�"�㓦�Ӧ�i�I�U�$ub���cH!MB�N&���ڶ1�|�4�l/���Iw�e�e�2ξӘ��� $@ۿgޡ^N]Pg�i��S���ظ�ކ�^��A��kt��h<�^�J���ZW�L���XΆ>���T���Α�h���	g���2��weC{c�7��6��s{�+"���&W�!���b�n���u1���#�����eU����j�EbG�s�ys��ͨ��<#E�)W�i��H�Y�a"s(��G~
���h�ir{~�9��MLf�@޶;��'�=E�'R��$�I�%�*���#��لa닙��S��!��<�=1T<�Pl7n��f[~l��;�z���Vma(DQe4[�2}����'���5W[؍�,��������:����˩�����T��G�s�9p��8����uZV��j�5{�����'W�u�+ֶ)��Կyd�7L��oG[W�w˰οoΜq�+M�2���|_�}� ��~~}/5f3l���ѹ}�z&��+�HtM�ɸ��W���#AZ�$o��^p1�O"�&�w��l2�~߱�Je�ɇd�&:�C-yB� ;C�/�N�H/��zEŞw�~���Ƙ�h�J�W�H;'����`��5��4�>�>���[�,�ٵ}~n��Zl&��{���>�1K.�&S9��0r"��
/�*���"��h2�:y�]#�J�0*o��E����#����kFU߽���S��Rb<��|ƾu��k�xFx�$Y��{8S�j�k�ʺg��٦P�3�{��|����� ���k~x]�r=�
C��{�eY�e�v��'=��ݥv�'� �ј9�7���M�? Z���U}��J�v<��BNE ���>��2�s/1��{�=�Ƀ�	�+� .�U�0�� �埀F3�spv�FΚR>`���Tu�ې��!��qm@���b,�l
�N�3�u��M <�5M���z����(�2�NE���Nz���vs�����y̓z�&
SAy�9�'UNT'��/���r��;�㳤sz�\ ���Uf��Ų,�ёӊ�NIQ��1���]3�ф;buz�Q�S�^+���h�w:�ZȘ���)Nu�����,(:DZ�צ�y��n#9S�!�c"�_�fϊ��G���wZ��c��
Zg۩�K�z9��9�_V��4��sOn>v�T'�10�����=����2���6���ƚ�!���?K�R���#ϭ����8��~�r���,�þ{�鱗�uů_����k�m��� ]����DnQ��552�icl�Kk��{XkS��R�X ��F�-8�Y��������}�,0!ӿ��C1j%�TBx)z��ݘݓ�|=�4�L>/��@�Gi�f���b4lJF�:�S'�1��&o��QW[�z��ւ�1IQV� ��yP�C��׀�Y4.�^��q�x�1���.�Y�s��i3S����7�`r������X�:�������X�Y�MX��yƵ�t�I�:7��6f�ߴʹIc̯<����>�Xj���|�p���C��hs�l}g�hdO9#ܦ��;i��<<{��'�0�RB����I���'.�q�P>#�r�1��p&f�+f�i��"�NyS0�2�����L���O�mi��!vC�ĴP�p
�3u8c�S�˲��M�e��*��'�������= <������N��9��e�(ul�V���Ґ�� �����8�#ίM�����X��EV�ݜÜ�z��d �N��z�)��v��}@;���������S�����zF�����|�s�Oy#�*�L.ي������&�~�:�En篏�Z����3kۙ��ϒF�4g徢��n��6�A ���E�r��6�����6&s�=����Gb�bf)M�(I!��s��, (���7��ױ�`���>"W�?ge�̐�{�>$O�@��sYQ�A+�������ַ�n����2q4H����������7��Ac2���C�~bDyٽz{���=���;�P�`he$f7�?�2�f�M��`8gE{N��ĳ����*��?������g�E�($[����U7���+!��`�:^?�x���;j��9d���o˛��9}��ќ�r�ks2��r{�!�L�1��fe%G���mx>��3��ʜa2��WH2B�Cv?�$(�.柜i��]D�6�������8�1P�q$-�)�|���ò��I8k6p���,ض�B����Y�=��-[�>�n�TG��~����!�l�I�=��ȗ|u��mi�k��R���BRڇС��s�D�r�d��|�,�3s�D�'H�v��n���`j-ge�<�-��z�f�m�I�t�\���X�d˙�[e6�PWm=s^����}vq�z�<z�h��Ϥ�$��{�3�5`����AE��#�R��������Y�t�Lq�����冯߾ׂͫ�Fnf Md�:Or���{m�߷�Ī�pU�Y�QJx�2�E�1��9م��Cs>\<�2�Է���Ǭl?��9kY��5�ڼ�7�w$�n�1�˔�7Ef������(���:�^M"�PT�}���6����/��ԅǘ5�sXo7�ŕk�Oዌ[��/xBl\��;}
_��1D`b�~�-�UT�fx�gUjlX���wM/u��he�Ȝ�G������{6Is6𬼑�n����i-=���8� �=�C7F*�#o��q�J��o�]����&Kj[z�9b�s�6{ �y0y�)�����y�̔g��>]3c�8��G`�*P�7mr#vUz�w��I��}ߦ����7�tLڹyB�~Y�ϟ}e��Vkw_�7Ɣ�!r�m�-u�5������ȯ��˨'��{d0S=�{�g�w�������Y����;��٘�L��~���2�d�����1�FX��?b��`�E�;�,n���#.qOI�1���������56{��Ŏ�Mu����lNu�y]��-h�#�����K�!�RO���롅�Lco���)�|[���̞̰kW�g�-�؝3�Q�3'�g���}}XT�\k�1����쉦�J�/���hv�O�q������qg�f>8��l^!GMʘM��m����2�ϊv���Ϗ�J�qOs�*Yd hs�W�Hi2���k��՘��C���hkE�R�ES9G�ӫ�ש�)_Q�+����M����=�4�@�#�X0������*y��?���7�2{���2�a��cwYk�c:��vÆ;�;�����9G
�2���	qE�>�.L�s�	����ሎ��g$���߶P:5o�O����ڽ����to��Y$�E*���]	z~E40>b�$�W�O���Wĳ�Q�j���Ö)i���[�����Lf@͵�t��+m!��G����6� gx�YY_e���O����+�d��*�}B{'W�o���T��s�}�o�VΡ|��+��w����s1Ɣ��jd���o�[�����eC�E2���kQF�[ޛ����i��J�&'c�8Xoٸ���������l�k��XP9���[@���'�@R{����rN��n��N?�� 6l��5+,j����eL.d�@:/�tԤ�A*; p��������;Wv��ʉ!¸�`�v�W��i�Al��8��rZj��Ea���v����um;�P(���s��2% 0M�uAnS�q��NxU�U2���UU�^�s��Z��"!�@���\d��$ׂ��m����0��f�9��5ՎK��϶���	��_y��R�b�5�8�m|�qGcص�����g5ڄ�	F�%�㤮�1Y�y�=�I���©1}����mcT� 뵃���e^����h�yb饶(��c9��\����z�I�iBi �p]u��� �	�g%���B��<����}i��^N�4�cr��=�޶m��~G��`��\z{�!�DMIZJ�`a̒B���k ��?`���A����> �}���������@{�ǈ�H�rk`�˞�����G)���3+�$k]k3��5@�A�O���i�i��P�ʞ���cP�
�{�Vqf��Q�(p���2�t��d̴ ��DOyo���G��&��y�@��?mq�AR٦���7Q�M��{�ǉ�"�b����ߪ�9P�*0zTF�Q�ܿ�kL�G%�n�h:������Ek��R�@�ٵ �6��u�2�Ƣ�Q���Ds<���yo4������:%��L�N�uh�%=��=R���U��es�ׁ^��+�q~��G�d�?M��,Kֲ�ݫ�GC���r���j&�s5v�����w���Lko�#j�" ��R=���º��q��~�5��.��p�6~?1F%<;
��Řfkܳ���Ù�|�#��<�Mu�x�;E��תּ��x�<Gz�S{�Lm霼{�;b�X׵�'�k]�,�]z( V:5�E�&-&���\�4�.@=�@���F"76#��@��e��j{m��Pf�c|���w.��O2Q���{�� ��nB�p��gy/CΥ���U��m؞i��խ1g�J� �6��9���1lΘI���!G�{�R�ј�sze�
=#3N��1N�<#!xDc`�I{�[�,C��.oS�j#��3�L)'c�����& �����F�%���I�R��3[��?F,��~��c��oJT~
Us�r�wx�S�,��&T{�Vhp�Q�U�]�,/{U\�+ye넕@G����t�'4i�$��1�����%gz��wv��ӽiﯷȼb����������$�bL��Gf	|1<��Ӓʍ�����y���G3��d��g!A�d{3�X0_�s�z�}�Fqyi�De�Dی�������y�rI���5��ֆ�ZuSo��lN�u�)@�ef7)#��TcRR2����}��i=��3���H��c�w����;�LB����(E% 2�����Sm�ny��������H�/,b���T�jYo�2�mU�e��41���hD���ۭ��KV�;�`Y�:�B(�i��<K�z��䏻[��v|Y�3�?��E~��Q�l���F��Z Ȕ#7�&Zub�����L�K���{nh� ������q�}�3;�ܲ­c�,��T�δ	8�o�7	��Ir�����G{Kp�C���.�Z��<uv�= �trSA��M�L�*�/��^M!�(n�qa���ܘ�s4� ���T�|$��sy.ow���\�;�X�\��cR��)����S9�y���#��A��B���h�р+��Č��C���Oj�s�Y4�mz�:�s�1��{�=>?7f�ls��j�fL(������{�����Bz�9"=_���[	��)�am��|���cR���{���.O�_���'����]�l���)�Od6���V��1&���"[tc�`.Ε�+��lKcz��\d|�z|fҹ�6��x�GpIByǏ��{8���m�yG�e�i2�Y�oۡ.	r�\��<ȩ�R�}�to1��Yg�z���*^�C2.��1F��I��A����6��j@��Y沖s\�΂9�s����r5�@�Y��O�,�m�c��F��g-M����nY�s'��<BΙg�j�;�|h��s���Q�;�c�k�ڜ��i!�,k]2���Wן^|��ywܟ{~���Ap��gÖs����1	2�����S�F��lNLV����!�!��.y��_�/�W������
���,?���ҋ�l�1��d�Y���E]���0��݇d��Ϭ0�vS,r��Lk�t5�<3�Dc.G�����)(�97|!��}T	��jZ@�N�h��Nʳv8g#g/�����g}�Q�P.F=�;���9�W޻�G�W3�g�E(�]��]�"�c����������lS��������ث�l|��Oj��B.�
.�~>��_J��u�Q�>����S�/�%H�u�*�!׳VSw�0y���`c|6�J5Ƙ�9�Guŏ�Z�?�H"!��b	��m�M����Rp@[l��et�LЂ�����������x�@! ֤pE��S��]O�GD�\���uź�t�����6wD�s[��aZ/��J���;�Y:���GrB���?�)��G*�����T0$<.�QrܗX��YF�A9Z�f��������f���+������su84�
�ʠ]Y�_��]ap�g�P��?��iv2{?����}�\X�{���W�E�7��n%�����Io׻��3� ��{������Hbs���T�g6E�FC�����=� �Q�m��w���&T���!$�Iy�oXAx��B���I�a�߭ˉg�q��i�d6�g5��m�q��|�Y}��d����<�h�@.����	Ь�Rl�H�AaȆ1  "b�;(%W�=�`>>��?,>n?���oR�bYW�n7$�E��3��æ �2H9d2�61#��co]���zpu���j�}��5X/�[2+�T�v�S|l�_�3BϚ~Ϥ���Z����^��RceҤ��S�W)�Z��D�X��c�s��l�̳k�s�
.{�J�et{�{v����,7d�&���(��~6�蛦cݼ<y1E@�;<So�1�koo�H�¨�*���A�癙x�\�zm=#َ�.#u8gK\eG��Ny�BC"J�q|�tr�O^c�9 ������Q�\�V�T��e)g}Y� H�)�WC�{�^M)(/��>�F� �����Z���_���} �	|�����	�_K�2Q�>���"�T�!�����'��z+�<�T�n����� ��~�����u�]�$ �,�u2����?�����:.p�>���k�5��Ӡ��G�����q�n�}�
7�vm�C��Z��Bhm;�q�o�a�m:cz�L>�h�Gp�<.��<�Տ)�2��~�Y�eK��l���ٮ���9\��~&o���ǵ�>�3}m���z��7�4`*�9�<�6T܆Qn���J��U��m��w������}�ħy�h�]�:u��6������p��@h����<�����Ԟׁ'�(_�}��m��Ͼc߶:�K��c����i�s �p�I����?�d ����7�e�� �f������gb���.y�3�J��0��d>�Pԓ�S��E�E����=ge�Hp�C%g.=�P����_�FR��g�h�`e6[U}�e�){�M��;]���	��*_��%����*2�\��W�ٙ���י/\E�h���uv}T�Ɛ<_c�s��({Y?�ր��Ͼ�Tv_Sp~m�S}��JOo�������m����?+i�icR_�dY�x���#���0��Ź�s��Ќ���'� �����,,�\�2��q��|�m����Vk`B�AXc��.��HƸ�e)�4����D�����f13lݙ�v�=�X����T ����d�D�l`�,K�F�8c��j�O���tt��ki�(�/�rB5�&��gsև�����&��U2{o���g'Yc�W�j�բ���bi�O���%}4�i�,��Tn��^ۮ���q�1%{��yϲ,������Y�>���)�Q=ܦ�M��lꉕ�u���������p�}?k��ָj2��k�Yl���x��~�j�]��9|Q�s��ط��~+�������ϔI5��&�X�}�X��-	�"�F.˲�ܡ@��X�=Ō��?>>���F�����v+;~���m3���D)��cD�pua��A�� ����VH�-ku��+�!�����^��\�Xk�vR�h<}L�)���<�e�=X�?�>8��6��IU+���gS^�>ӳ?>�3@����EV�3��@&���n�F���ź�7���޽Յ�%��yH�)ߝ�3g�S�L�g�]{�f�7������d|L��=�(��M,����5�q��S�3��A�f.Dj��M0���3i�x[��~OW�gi��W������X���Z��G;d'�k-\6��u�!�b�G�T����;FI���W~���l琘�������{��H*��XZS�0=��2�[�R-ob����G�<L�9��R�S�f�?z'��]���d�?O���eN-Z'J-��5�6�V��ڜG68�g�t�`�����r$zh�# � ��Bi �Εj(���u*N���靧�R��&#�h�HF�>#=`"��j�Fn�x�i�Ec�^�u�̻��޽3Fe�q|����JU�����ˆ޹c���=٫h71�^F��:�I�G@/�S�6s���cg"�{JauZ'C�wz�d$��Y�������+���}�ض=��M�^pE�,ek�����_�2v�K��G�%Sᨬwɛ�خ)��ɀv�.�]�<�� �������#MlLrPRD�l���v#[��r���^�[&�'�Gd�Fh�x�qt*3��&���l'�ת�$p��z�VF��p� �jAl[/�<|T�#�DN���G������x�G��-B`ʶ���'�'���ǆ��)�J��Gc�w���p�]ί��6���<��zVR@&W��>?ڿ5��A��G��g��X�X<Yg��u �xBa˾�OP�T'I�(:�8�e˺����%�mm�6�PB^���6���܏������nQ����%� ���A4�`.?��=��K�S����� r�K�1v˨;>)�1�^-W'mBz��^V�Ŗ:������>��Ot!Xx��z5O�6��=]��bwƺr�E�qƈh�Ve,t��|O�ԛZ�U��g�e:�'��3;[��~��9��=y����s�z����/���r�50�2��RJ�ׁ�B?���6�wN8��A�������U_2�� I���x�1����HxT��F][���jG��nr~%[̳\�=��4����}�RD�;6��f�q536�M�d^�^4��&�����v�3��������I���"Ę��1�cROJ�f�!�	1�܁�A�#<�q��)��� bZ�mD��zĸ&�-�b��G�88�L�~rg�^cT��)�Ĺ] p��w���_�;X�1_�E�B��I�v�1��������Ǐ�#��m���t���I�=b45N��yā�bz���*�x���^h����nq9[���ю��oe�Z�{m��4��k��ڢ7����1��}�����<)zE}5�aUS�6��=���<����j�to�,��$5�y�1�g��ʻ���j��1<�z	4��D���s��~��	�T&��Ӵ�V֙����c�r�s<���1NML�FD�]wt��$�3R	�Vs4�s{e��?2��z�1	��)�-�q�L="|Y�,������m��w��l�����<T&3�����+_.o�!���`��0,4D!���2���Ao��ؽG1ن2�1&y��Ђ4�;��su�8m�����@��[��'��ф+�*m+	�R����=�c��������LNz�����W��Uр�"7G��ӵ�-��$ṕ���o�~t�����ض{��&#	�YP�0zr�1�g��d���>����)���t��^�)�y�{�&�lm�Mx��Y9���kc�7�_ap�<��
v��_���	�g�8����/ɬ-�\�$�;H�/� �q'�f,�j��)1��O������g� ک�x࣢��!'�h>_�9 �mK�?��q[o�9���kq���I$��M��n�l������v��)'����y��f��1�l�H4o���T�;Rp�7)�yP���d��M/O� 9���Z���OB�8�3�[��YPp`��v�l�_f��w��l%��=��9ڹ\�w-�q�S�S
j��5�3cL���קd�d�\���Ǭ��m^$�/�nۛذq��J{��@�gN��C��&�����h:�0��8)��1�fY�0���Q�ʌ{��\�-SK�ȼB���h��|>����e��k:K*�9=��o�1�2??�������M�9�9���Jz��8��YM>�����V!	hR3���ʹ"G6���O������#ŵ����UYǐH�e��,#�1Eܦ���e�!y�lM)���F�e�9I��m>y��@����K�;����\d���!����o�Gh�l���M�d��{��/�Z�UZ����ǌhb�a���H	3���|��8�Ƨv>={:ަN�B�}�M��5ᠾG��o�}Ed���*���
I�`c�d?��v!���0�SIj�m�r����v�aYW��<w�呍{=�ډ��k�n�uB@���2��[@����/cm��&� ��6&�CD���ù>&�K��r�0C$Ƙ�c��-61F,˒B&�A�m�����z���TˎD�}�S�k���u��4����nXb���#�T#f��<-t�H�%��Η^�����E3�#��M*��vk�ʚȺ5�s�ğ�/o�M�m� ޳�j��:�=���+��#V�D�k�]g�龩�uu���{'��#���8s0/��� ����-�;����@�+� ��?k��w�[�����5���-E鱘�I �=�+�C�N� Һjc��7�}̙�%r�Ǐ��~/� )����a��{D�y����w>�-�cL��t����\׵�1�([z���a�g#��������s�G\\�Q�Bܷ;Vk|z�>��>F��)�j]UdW79v���(�1b��v��ݜ�Uzy�-����T>��uo`���h���H{�� �\�s̈́��Iky�eZԙwq�f��ې\�c溙{���Eq�c���h_��/��?�j�*[2M��^�+.���F���IjS�A���|��z��B(���{z��� ��J�Mb5#�c2i�9>�W͝�!2s��"�s�B8��CH*�I�U��h�gbg�&��o>kzJ׀�WH�/zH��.3��K�_0�G��uر/�"�Ě���- ������uJ�� 4I�gD`2Ā��p�|4%`z� 3�lL~�|�&���B�9�\+�����Y�`Ɲ7ƀ���a�w�G�+glT�sի�Im:f}�*�dS8�1^${�9ںc�K)ŀs�9��H0�Gg@s��;k�3g����gE�w~�2���t�
�_�����e��pUm:G�W�r����y&tg �+��L�9
���"f��D{�[ۘkeʹ3����BK������H#³���|w�k�Jd�w)=�)Ͽ
H���e5��:�>3>5��c��Pr�mzΙ���@�M���}�~��1"� ��w�[�2��������iDH01��(�YMxDĐw1@�Ycr����K�!{�ֳ<�3�D1�/�R�ҋw8#Z��WH�Qm������z_�������Β��՞w��ب^�]���^��ȅ�{K�{T��u�rfD���9Wʓ�������7�3)��w_�@F��6�^9�lZT�>���3o�^�G��=��ؕ�w�3sy��>&��E�/7jr���W	XG��-��.r�@qSe[zk��&����xyd�ޛ[��N����8����&��5���U�Yߌ$O����寔���=k�&#&Dk`qd-�۞Yx*/���d-Ƅs�w�[@���������KU���1-�B�-C�����n�ۆ??����l�3Yif�`�*T�1)��8N'��1�����>RG�xg��Hu��mr��;�^��-|Pq <����1���ߪ)�zyoe�u $���e���sIz*#�^���:���2W�s�M�WB��ލ�.������� d�y�r����???��L����dy��BjcA��[����8	!�vkճ�W�#�l]���_��Z��1դv_uө35=��oV���ۆ�x�?z�{ M���ׯ_X��8��9W7��^t�oN{��ӄ"�6£�E=���^:�w�چ��m;��܈�́����oJ�I��)3M�T
U�	)
uQ8��;� �y�u����6t�̝H�}ȱ�˰����^�:�"�uŶmEM�,KJ%�m��ׯӲ�L��z�k����c#i��|�WvF��C�2����������_%�]��oң�L�����vA�Р�`v���ۿ^W��DN��:+���,��h��ڐ�imiZ�0vT���Q!6�9�u��`S�����1R[qvB.V!�Cn��&Ø��M�۶A.t���L����6C���7�j��+�PZ���b���_C�#����:J@*��}�5Z�l�����.Y������{�6ꓲm��f�ߙ� ����ɕ�]���ujjG�V��HʲǦ9�&���c6�X"�YY��O���sh#Z�Q?c�v/GR�:h��f���8簮K��b����XD?!bkPWs����uY��;B�>{���j��w�{2��0�X�X�S2�� �bN�b#z D�7�s�۝l��r*�� <��X:�l��w������F£қ�_�fXO�5Sl�t�ƭ�ؑ���n���ƺ�Z-�9�c�{ ��yZ[�B���ϣ�g��e�">�&�ْ^}grD��͐&�j�p�.y��H��WcO���p��eaX�y�ڔi�L�/��1�4L�,�������j��K2��5��Y�!�*+��y5��(��d0�
/����]<0ۓ�T�&Vq�n�=s�Uı)�U)$g��W�%Ùkӆ�rn���	t�y����	��u������Ȟ�(z��K�=_bQ�7GlmNH{�/�9�.Tv�:�&�C�a����}?J	��%ˬ���蜅��0P������pf$�{_#�:.���A�k����R�=roMFޟg��>SlEΜ%u�����!����0���J{{��^9ZF�l��]��P��J۶I�nfA9kw�=����dd�^-��^���U�d�L�h�M�T�4,���`9��X�d6gL?ZV���>�,�n��Q�}����~t��DS�k��.��ym�Q+)70Wת�{���i$�{l۞W�p����d�im��ub� �HP��X���L�# ���1Tv1ƈ�}
�.���Y �K�06y\�gN��̽�����? n�ٹ��P�!9�P+�uI��T��xo�T%_�t\[����;�|��׶<���7[ՍTy �DM;bT��k}N�̄<�JӤe�P26ݙÓ�b'a.�F >>>�	�"Ͽ#��(����j3�i���V�<��m������y���h��������]�hA�e~~�Rd=4'�M�X�I���+��z�������L��]���<i������]������Dۜ���m���9)1���[Uk��v�TA
%�H���V#D�E>����PW/�GO��)e�����\��_�?���"�=I��mC>��\�&�Z�b�v�b�����X���z��䫂�I���L`�l��&��&���E&A��Un�a�~�m�v�`�'��
�b�HB��@��tT���8��y��r�z���2A��,��v\����-���#����z���Zkؠ�ڽ)^�5��o&�WH]0hJY���\z����CqfQ�)0�1�^�L�'����Nm#2f�̳w����Z����~��k�P�D�(�|.<Ǵ���e�_��4�����Fa�~Z��=���W0h�1�Y��d���ό�o˹� C�	�P���YR���������ڤ�F��q4��:#ں���h^mLd�s%�9R�X�\��q_�\�٤�w�j��g��|DM2St��DI	p��@��8� �J����{l2,K�"A�9)8{�1&���mط֤��!xx
-S�� *��p#�ir��9�b�?�v�▮w��6SY_:� /)4��fUL�r�ұ��o$��%�Ag9ؒm�;��}Iu���]f/H������#=ïQQ�0��-r� 6Ml-ȥs%c�7bG��'�t��}L2DԮ��F�� �6W#�X��~����y�{�Z���G���T��%��ff0��j��� �:���Θ�̅g�c9ɼ%i�b�nQ�5�����.����p��ކט�	7G� 3��T��Y���a>~���?��ր%�����,�L��献�]e_�~#�Q"GR?��iͷ9�����i�N�8�يǫ�6�r�H���u�PC�?1$ ����n�>&���@2�){y�	��=E�wKB�9)2F����r~�ٞbYWXWӒ�vɩ�&�(�m��<|eb	���A�c�fH�N�r">.���ec�����g��ԓ�eU}ulǸ��IL�Z8�c��d�q��Ť&�������i"'♸�RF�5��c���()����g%�5b/g6�(�cs�Fߑ
7۹vOUe�,<L����s����~S'Ǎ��M��1��T���q���r5��Xa;?�u��i�j?9���(c�9��#���ػ���;���s�������W����v���cJĎ��
%����[��9]תt�)`|��(� Q���&o��,v�q>��f�`q�rg�sn��9��β�X���0� �T ���;c��������vq�Y����c1Θ's]�!�� �#H>.�9�69�1"g`��y���0�I�0H���s�׎7 �oRQ����9Z�8�*�i������/�t���|r��uml�t��?�{F���s\р�y�\�s�1l�i �瞞]k�Z���kX��9�xd[�L�Ǚ�^�99I�T}�;-V����T���&y�Y�n?�=�9P�1�#�Γ�;��0�A���{��:���vks�L��랃��\�|2�3c\�lT��I9�,��`M�������g�yI��~B����9m>�[kK_m�!�C��m�}�e6�|%�1��X���?�E���գ)�נY||| ج��=lvh�sRm�������1����{���ᢝ�w�{@�������9$�S�	�&�W����-���/||� �:9/7��`��ރ4���
c��Eh���R�t�MH��ψh,����sz�=ϔ�[��i�&�����3�����˄�}@��y��d�S�Eq/w�9�m��W����g-u����k�ߣņ�M����#�N���˯h-`��7��8;WJZ,G���=+klI�f3rޒȾ�5����إv�Է����k{���Q$	���8�HGyUڍ���FK�栗w�����e7��+DK5y��$�;݃^���q�<�K�o�ֱ��C���9#BF�!3����~���'���w��y�;�୅�d:�^H���9����!�P@& �l�@��z��D��������O�>�h�����!F�9Nf�X`<�8�tn|<?��A6{�#��/�3��g�L�su��-_g�[��M�q��R��Mׇ�S@oq�m��g�&gj��vj��z�^�S��{1�<�����q���<�ը
��U ������7��֡���c�g�~���@e��@�,(<��-#I��WH��5����K��m�!f��+ޭ�Z'��fϬ]#�r�~�u��.<����s�q��!h4>�I��s��'$&��^]�^��|�ߓY!e����!���	�:*3�_Y̨ ��p����~/e���A�ɰ�wL�qc�� ��6�'k�����Uy�)-$r��*���9�Y����穩x4��i�z�KMd��z]�Kg2
]�Ղ���F���-�h�-RmN�0�ɟE���@�4:/e�8:��ܦ��ۆ�����*p��^�*�?^�,r�TOzF�&�P����3
at���^�)���\i3�ִ��k��P���@t4GM�ݳ�V�Iɔ^}n����߼�z[��}���v˸?��g�u����xt�����Z)�L��Mf+)���6��j�2����&�}��=���^�i ���!�坖:�.�����vK��� ����Y9|�p�U�i�^�4�T;&I�l���#�������������'~��kІ�ޑJ�х�h\�?�H^����������������La�\?��#��l��O�ږ��m���E3�P���t5���X}W�x�ئ�Q��:_=�֞�'�7�L�����c`<����A���;�d���G���Ve�2VlO����<45�pr|̜�������>�!1�A<}\I/�U�mt���u�h�X�@��-K��U�i74~���Y�ڔg-n�[m��܅ f,b���ܷ�X�e�-���6�˭E��a��pD v'���;~����!�c���c(/���@N�N ��!e��[�ݺ�X�������nF������ym{���{����QF��S,2 9���t���+�� !@޿�!��|��������s�����)���~#���h�!h~3S|��D��H�J!I�1��N�i�cU�ߏ6�
&��I���t����h��:0�·M	8H��B9�p�J�����^ߔ�'��G��7;o�&���g�}����3v�'���r{L�l�<&%�L�d�Fʜo�^�K�;�U��NMDJL�t�xX�v����)��?Afcm�n�10�v�I�@�����p��:h�=b��!�f�8��䁕��)ʤ�{lv��v;��6-�$}~u@�+Ҫ�	@=6g<���gκh�/G"C��������z�����ha����jR�Μ�#C�k�t@��΀�G��2���L]�2��,�d���2��Idv�ٽRx�@�����x����c����1F5��,h�x��n���~�p��}?e�ly_%\��L@זѵ�)f���`l�kOZ���}h=���t��|����@�))L{�T�dWIuQ�6��.93�yn�@���ɛ��l3�8�����0�M���)b��c<|��@�]"2}������yJ�BL;˼{S'�ض-��5�dv����Z��;bf4��u^�K�:�9���$Ay�[��\��
P���_�
�\�r�>����j{m{����WA����Ũ�����|�	���71��lCF�EPz4���X��ј�m�1���h�I}���5u�loe�b�u5@�dйǯ6�zҏ�aϏl��43I/�e����ȹ����\r6�iL��z#�# k=�9q��J�r��>�9�����;i#aKݼ�kz���9�3���?)2����OA��ែ9aM֊�
�c�5G,���"�� =Ţ2!�A�3!��Ie�^
B@�9Ŀ�Z��rn�1>�ǌ1�mn�b��o\�񷟸}|`Y�#���������Ͽ!�ڔ����V�[l�ݠGv��2 �:oo�׮��ˉ��m{�W�F��=�|z�6��O�`e���N=�Fvhb=ډr��0�T�#�:�#�ʅ��h���l2���c����6�#�X:	8p�����P�=*M���9������ϟþo��O��M�I�?�����~��\�Xڥ�����1f�,���XsT<nRS]εv�������:ڒ7;m�?΃�s���lԮ�ߞ�0g�2{D�uM�l���\#���@���g��KnL����G�ѓ̦,K�9-iQ7#Ǩ	L3glb
��[���5���sr��}�[\V[��}H1��m+�ŀ������b]����������}�@BL�g�/9;������?e�R.�f��bX�O
Vk2w���h��SL�`, �)m�D�8��.�R:�lR���◐��H��Y�t*�բx�Hh�]i��(�@p�X�N��K/�3y��\g2���D�t�3�[ӂ��M�U��!�D�K�k<^g{{@@o#�M���r��ƃ���5쥬��� ߋ�X��T���3g�TNk�Jy���Wz��c Ƴei�i��x �c���H�F��՞�t�y�h ���M}=R�|�����jWZ�BNf�u�e5Sl`J�x��n�p0�⛞ѽP	μ��Z֛�SO$�X7�IM�w�w���A�61��'����۞��@�2-��|H�7� �d&1 ��c
�l^mDy9��1l~�5���Fg��$�Pj�L)t<��`2�or�{|t���ͨv�����:�ɵ��W�[�c�?=�����Q�7#Z�)5dR�˖�s̳jH����#*}�jH������PET>�pkZ���ZAΨ����<��dx�g9�]/ߣT�ҳ�D��-\ͭ�k��S@z*�6?��v��m�@��繻�\u�Ѥ��|N�
ဌ���W�ن�;]>#��	��|ޣ��|<P{�1�M��
�v��Y�`]L��ͻ��!A�F���m���_�����!9���?��9�xDާ.��������O��D����Φ�&2� �=kw�Mgg[���,^[L�DƘd�˘'�[��Rf�	�ؑ�H��h�8��H&�jg�X���W��Q��홷��e�ꡖ�!O^y������V�y����8�@�
��HO�I�R�5�}o�Y'���1~�HWK!����U�ͱ�|!�߼,Y޶mͱ^����=��@S���9�S��ϥ���A�3��y�w�(��T���|#��Z��JU��Ȁ���; i���Ƒ@!7}�]��ly�@\��Bkb 7j�Y��w�3iyVl�&����-�����G��o�²��.C��۷i��h#���d�c����Bޫ.�y'@Xr����43mR�X���jW��-�7X��^P\�߫s���>�}�������>�0�ۊ%�ق�a��� b3ir�~̑����F�_�b�ߥ�E5�'Ğ���T��<_.�ς>	���Sk��v�>�̲��Y򺠷*�V�Vw�5/|jǱ.��m�E���$�%U��5_�=\Oeh�	��CrQ!0��J�NmZrީ�Z��{��!�ڮ^��h�I��/5�K��(�8/W�;�C�CG�pW����瞿�MzNM8c����T��Y�s�5��jw�e��`Y��ҳY�NË��Q_��9CO�8j���3��\�%`�v,˱�pf���i�h=�S�s�{降�k��MM���Z�m���0E���%���-��c7�Ԏ\��X�
;��i/�۶5��i�s�U�m�^C�=���JyoƟ���<�:�$����zM�91��[�X���۾cY����v�#v�c+�uA��Pf�y�
��"l'L�� <�����>�y�C^a���J9{~�F�����_���Y�Ŋ[����B]�~�&;Qk��9z��|����=���-������c�x�>8��3���o6������A�8�Houn~ ��z�\��j8*����Y�>*��|L�8���{���6sq���UB}g��S{���s��{{,v��6��������6$HԀc;gQt�10 ��s��Ew;֤2O�͖2�hm�rn��Փ��$<�m)U$�Ĭ6'�8�������o�ɴi�MJ6�Df���DĘvч��˨�Yk��;�x�|~Q1D�o;���}r� ���h�+����6H���˖�E��N2i�8����
�ʙ�������s�W]++s�����ZF�;M������|d��qN[�[������6�>O��4��'���T�B�qƦ�3��:��  '�9���]|����%�n��3��s'��Q6����Y[?S(%�!����`�1��y��|Ł��m�;�=�L�l�θ�R��D[��͟� i[B^O���eYA�]^o_�}�m�e���l�{'���Qנt����-%��}K���{)w���o˼�'B�@�(�zb4��20���߰�_���˝sp�"����Dǌ�?� Q� ��4յ:��u�[*1���E�a�#s���=��*�c�Z5��=��(98��A�[F�W�G�Z.gvKg�>X��I������IF��G�yVZg�
���z�e1P�M�����G3�s�є����ʾ���98�$f����N	��8�,۬��������H��{���˶��,�;�kd�����$��z�S�R��Q��w��ߚ:Y{�u�R�LT��,��c���e��}ӳ_���Ek��u�m��x9�y4o�֒������q^���9E��-K6Scjr^N��Y!6ӹ9Sap��Mb��Qx��6���$Ǟ�h����O$R,���;d�͎?6��<��$��t'2�u�LeF�Ӊ���5�q���I^w�{l����cvR�~�����l�����D0䏏�Xc���FY�*3��%#4���P	���rt���I�׌��m��J`2R�h���w���Ȥ�s�y�w=u�Tk���z�؈T�=ன$���P�>�?��|È��jϹ���L����;��:�ɶ�����JǬz}�2�@���o�xCժ���Ӏh��l�ϕ��*�=?���9���g���N��e[4�9�H��eq��}s,��6�Zݳ�������@���b��+��ze�R%Ɍ#�^׵�',}��0$�~�71���M
�,��t�l>��!����a�n�m�Tv�������_�|k��9�g`�rb��<��x�q[o0�b�q/��%1���, 7��7��e��<������0���LOG����P#Q�Xh��� O��rc�tK��&�~� s�5�� �)��Tj��XG#�k P�t�ݪ<4)Έ���G���M���jj�Z�װ�='��.4�p7Է�5=��3Y5����&m�Z�u��[�E���g�e��|y���>sxN\�zt&��2�$_�[��Erg�́���7
��Tp����w4�0�����^y�ʛ{ɶŔ��5eh"�%��~��m�N�h���,�Wh�X�Fhx&����-x�˔�is�,G��;����mrf�,*����k�a'8mZRmgB�����Y} �پm���8��?=W�[�e���;�ƨ���2��`����yƕ�0�Ê8��r��*��$�^�:���5�j�yd����# ���c>+��;>+gf���'�A��=�:3��"Ɓ&-�	z�|8pЙ/b.��NT)#�����k�+�2fG�A���;J�s�����)�tn��/3�T�|1� 5zv��!��Qbb��NK��7�5B��9�8��ro#+�����u����b��u�\�����5���Ap�Ϗ~=����1^�������3�C?�$2�Y���\��Y�=�>���k�)��$ۂXaeb"`�q+睂��$C@4&��1B.���a�7�=e�������KU��IAg�����{�� �����Q�N�Ѥ ��;S���V�ދ���1����S�])���
�3_c�.�G���v��d53�����衔�#���I?��Ř���������M�Y?���ҋ� ͣ��U�������we��X�u�W�,��s[J��Ȑ�{��`����ׯ_d�W�7�3"�6���B$��6��Go_h�8ק��o�`�[ǌi�ͷ������s�BϜ;���4q�:�N�>����ڒ���cyZ�Hz�q6�@��>�56����\�2A�<�$dnL:fR�t�����(&S�d�cDP�<�ĺ��yg0���Ǐ���'�s���Y,n��v+�c����b�5	�z��s�� �@��I�7�x(���gw��$,'���I��k����~hs2�n�6��a=�({ A�П�E[�Wp�GK��z@C2A���3��gl7@�f�Z\EY��MR��5&�����g�]/dO���I aΆW
g�y��!����u������i�wҙfdüm#�����V���1��-m�u���������/�]�1Q�h��q ���C�6�g��-7���t�S�x	͹�޳�,-.+P����b�M��@�$?���s��cYֆ����~'�� g����H���g�w#���}H�m�������J��(g�q.�|4��:cL�rc�Lb"���PF��5��aM�6�v�H�XlL鰨�`bR���w4ȕ�u���Y�}P#W�� =��+e�<c({�H��US>�9Y=q[����jէ���{&3�L�=z��E���I�����Hd��<��;2?�67��a�:�h�9s|� �>���6%��3��Y�гe���+�Ң��n��i����^��I;r	Gi|��kHڌi���v�P2g�7�Ĝ]I��7�Z��(����k'������Ȕߍ6���+�L�5Ҋ z?z-�y�!�CS	�4����ڀ�G��,��7lۆ?���9�l2���%o
a�~����Xfc�����D�}�
���2'����&9��=z��|@��to|���RF�I���}0��;8�o9�[���.�Q���������W�>	���b�O�Ln��=��M��7>q��N��,�)�|���L�߯eo�C%q�A��|>�w�4�cc2�0A�y�<���*��q�������=e�y��t����T˲3�/�����[�c�K�s9��o���K���3#��w�L[4�����¯�ŕ��D��gs��I�d
��=�τ0�1��=1�䐋��X�ۯό[|�����}6�Y]�8��Z$ԙw�����ff4a�r��#��i�JX$c�
2�ISQ4�[g�L��v���v�\x�5RYs���(��������~83y�M:$rpK��,CSm�/��U�)���¾�v�J�z ����uÁ��#�3��K�He�jve>4K߁�������xp�����[۲����e����g���}�j4i�9�ݮy�˺�߳Ϙ�A��G��h������;md�6i#/|�=�ƍ?�Q0l�	��z�|�o��B�,K�"y1�ǣ���J��2�W�Om���W���+��J2�zP�^[F�͆�Y���M��yDlag�_W��|)�w��� =����)�4|���w���)��6G�q��� ���1���Ø�e1�� ��˘�&��.+ֵ}�����|����eM������vº��$��ý���XPP�������#�F���$�k���F*���ϴGVG�L�l��I�+�٩�́1/c����+��g|��Oe���z�f�X֚:{�w��P>:�>`�� ����:jʧ�<���u���G���9�&PB
������q�'�6�RF�	�s�z_r��_���y��/�!�CX��B'#�]��<�ڪ�'9�g�i�l'�}�¾
�F�(P�R������˟�1��$j��ևv��ː�7>��9YqjL�,�؍n�,˲b]<n���VJ���ƺ1��
ᅏ����H�#O�h'>??�g��k��;6H����d<#oK+�X��^�3(��	@Lf�Y,LLnB��m�q���)qV�n���m�[�c����u�*˵Ϊ�C4h�����BeK�R�I���BxFz�Sl���O�=���SކYV��g~L��Q<�4A����M�u�Sy/g������������<��9g :@�ϴ����v�&����+1J�}��e���'u�F�!�a�%��XZ ɼ��9��~ִ�+��鳛F��Ѵ'���5W�8��z,��OrК <��g�9Կ�10������� �>���7R����)͗b�`�RV���Mǁ�ر׵�?� �@}R���̘Ҫbp�����F3���d����_)s�!�Y�8�@���a)]�����
M�~O��&M�v�1��mn�-)�ҵ\�',>P@����2�����&/	"%�$�pV�d<�� �Ǒ{��܈������a{���?*�v������B�3��u�����������;{hʶ��A��r?�*��U���g3[��x�?s��Nyt�4�o�pV�
�9��4mǣ���{�����<�j��}�$���hj4߆s�v�,bt�.$'c�B,!ı�O��R<�RB���e��g�*��e@���>}~�_�A�2C�6Ĝ�'��={�ـ�.#ZZ��Y�:��[R
�e)��YDRg�y�b "�"1��"�;Ӛ9�9���.���3��A�UJ�����'�]��wG�-P��1�r2j�#s��p8�J��q^�w�TW�kW�}-���3���D6��A���Ui�n9S���g�q.-*�T�c�*1�pR��q�M����.�����x�u���J�����?n4�4P��EӚ�u��l��g��G֊g����k�w~��ԉ��}��bT�(�}"������rkUaR;��k#o���Z3y�r.$_�F�L� �o%��Q�l23J!�ƈ��!qzA�#�l;Zp���Ef�ͦ��,��[W�e-@����0;�uY��Ͼ�)]��n)�?�Qp���NJW�c�"J����� �!��Ο�f�$�#���1�wߨPd�3`X����|q�a��y��K3b�t��s�I[��Wdv�?.j����G*��z��c��k�3�ˬV���L�o	�f��ee��o��$�����I������!�������.�1۷����v<������I���x��aĨ���c��I:�0 bY�����u��7�bL5�~�&��:Ւ�* RC��k�oȹ�C�}A��}� ���ͳ,�񑄡s���%GS6�L������ R�p��1��~�= 3°@�)6e�l�`�MGHf�Tȥc��
1���ЀTMF�	��8l]�6��B#5���g�E<{N|`[�?n+��lw��&�޳��h��->|N��SN�ra-�Dj@Qk��GJg��WM���x��GE�����_g�?�]�X6�Ҿ"�ϒCBOz�� k �lO�SZx2�!B3��su�\h5�4�|i�������Z�O��c�N %�+�������0:F��Xf�Λ�����0��	��d���J��7���3������_����1�T�����a���~o���zy������e6���J6�R��7d�o�!��>��M`a� �q������7��y�{DĐ���:�Yk�<��g�:BP�L*bL�V�߆�0@��y�`Ӌ��C\�,c����	W����ȫ O�E��8�5��4��YP��3�W�G��&��޳}�>�̀���0g�f�Y�6��������r��רX��q�*���؛��8��$���|���{J���M��~f!���F��Uv-��!9N��P5���.��� �����A�	��	�d� �,	�e|_��~zq#{`�+7��}$�� 5P�r�i��?6�5@<��4N�>� j����kSGu ��� 5j?!����7����u�U�6u�m]����`u{b
F	��i,���:2����5���\���}& R���1�d�P쯖����F`��K62��r=�ց:y�v�i�7��� ��7ty�2~o=���Hm�M��J����W��D�[bd{g۩-��w�3t�|&��f��L��+�"VT�k���h�\c�����zc3����,8�Q}K@u���P�L9>����G���Q5걶��{�eis�~��B���j.ss��f?��q����Q�Gυ&���kY��u����� `i��9X��_`����|�Jzf����ߗʺ�6E~�y��{����ۘL#@\@U����%�ز�(�A����򑘱��z�auK����#�;��ǿ�뿦\��#����-)���v+�g�i!lt�`ja;μi{�G h'!�i��r�_�����Y9��1ǅ,- ���7�tk+6�2�sϞ����j�@��kc�֓c��S�I��Gl*y����~�E��<o�h��_�@Rl�6^�qJ��z|��# �e�g;���~,��1�n��M�4`X�h3F��em�i������M��ۚ�8犇0�ÙA^ߨ�z5���y�k��J�m^�k	�;�����2��=gMF�N~�k�d(�����>�ؤϽ9��c���RF����4BZ���1�ei�*kbx֘�.���C�ߝ"��=�#� T���'�mO&~��C?̧��'�����U�1���Y��˃e$a�eĜO|Nv�����g-�eAp벦���u]���	g�TNn��+��D��eq�^�L8k���DR'��ȃ��	��뱦r�Հ��hz�������U�m�b|�P��3�*G�ʶU�ʺr`1��������*�/sI2(��3I����=2u��קk�l|�c��Cb�I���w��N�����s?��iv�]����}DN#��j���̼}֖�hj�c�s%��7��}��^���������w�?��H~U��6<1e�����'��a�@��ӹ������=LfDyx �}A~6$�sθdp�ə��E��3i��=��z����|��er�g�9���b�K\�Oo��G�(Was��Dc7��Tc�4���Z�c���*b�٩'���%���^���3+�nc3e���l�\�u"P�J9�Y��Yc��ٗ�<��k���#�x,tN�����<����wH�mR��Vם<?�T�g��{�[[�.g棳�K&{Xg��wK;�s��*�
��q-��8��$��Y�%7x
Tֲp��?��:=K������s����W�9~����Ɍ��DE�lȚ:�CD�Ki`M �M��"T;� ng��і�Z2��,K	�n�Ų8�n)�:�����R����Gn;J6 ���O&��ī-vgO -,���4vQ~�TNJ�E��쵍�n�LGR�3��]S=�D2���gTN\�h�p�&�G�0P����1�ϲ��:�z�sPKm��y����9H�v��5mxV�3���1Vr2!hMXf�l���z��y��I�yI�72{�~;\S4[���f�8�$o���e�����ٹ�n��ה�B�Nc$U��S�*��^�H
21@�c��L�v LV�������I���������{f;c�#�,�&&3OdЅ������d(���I���)�޷ȝ���q[o���Ǿ��i����g�!�{ �_)����$�b�ӄ���M4Z��6�Z��i�X�n���Uk�:�!�?�xoB��/��~�#Дj�c��,�G�}88͌��u;�p�}�7M8N���y��~�ޯ��Q���'ߐȾ���,O�_O�~e�	��%瑞�͖o�ƚ�B���������d���3X�|~~v���j������g��m���Gټ%�z�����_�m���{s�6�̴_�{n3�s��N�W꜕Qy�1��[�u��1`N��ٞ3� )rL��d�x6�c�`R�Mc�S�j�+�����-X֥�]�M��w�d�g��yvT�1b�{�/d�S���J�f�B�! �����IF_�E�ɾ+hA�Y�xP��K2���06�ƿj�l���3�R]�]J�#z����c�	~�V��7SVO=���^+�p\Hϟ/�
;�
���I�q&4N��x��^���#`;����<{i����4���A�:��dC�d��x2;�Q�Rf7����@���ʻ�1�#��wچ� ��і �y��K�+kG��q�ρ�M��W�r�	@q���Ϭh�	�����N6���Y簸��pý�������fy�MfB��'�w���1"�d�
�<9�0�u�/Ƣܶ�-01�����5u�����Ӑ^���j'�!���_�|�3FN�[������l��2���9�g��y8W�H��w�gۥ�_ͪ缢o��2##U��s�[zc�����PbW���b�
��&t���H�G��j^!��^}) ��\AdĬ<2�xD2S���M�-s*��g֥G�y����]�Wu��ӽo[��:��~r��L_z�T��_(�7����k �{~��#Lj�����%��nK:;"���q)8j�\_U��z^3	��K*ɺ�%�芽M&��E�19��qOM���}i����Fy���kl��`h�r�}8c^�����2�W�Q��3��̵��ɬ�N/�_'��7�l�d�a��5^O#s���vlۆ?~��J��#re u��׏@����6\F,���R�|��K���:4�9��F����X�{_�p���!�F��?��bvLNd��EsܵLf{�}�ق�����!R��۶U���T�'�痈�V2���`PT��<��0�X�)�;�c�� �Rm��u�)�h�v�q������V����s�������
��n� �%?�c��\\i�ZY��O���0��+�&#�Z�$	Զ���"� 鸵���iǫy�'�L��mv�R�D��kG�@�S=�j�W,�ia�9���(3��,���^������:�C�&U��P~V>?����Nޓh�m��犫}���އ�v`�a�z�.g���ۨ��:>��ZgE�m���}||L���Y�3D���s�Ų�jߓ`�7fe{�9��)��3��kF�u����[sA{�з���5폼����8���Oi�#����u]p�������mǯ_u<n�c�6���0���1`]?���%���6#�SmD�ED,�*�޷��#x�",�*��e�3�b*+3HO��P���Y��w!YK̤���2��5�h��yq�k���̎R�9sIޡ�?��vǖ]i��9��\{����:�!q4\���q%�B�$�Q�~�Z�j�m~������Q�fh��sU������O|m�6�QZYrd����s�Q�H�5[�)�У*h���>�!�:�Z ��Ʀ��L�In(G�U�1+�l9�`2?"W���r�c0aݳ*3�p��h�<ٖ3מſ7L�Y�?�|U��5�|\GKf���*�I�Ù��a�il,rb�̳� �~�o���?s��r��x�0��x����������yg+i���CS�U��$LJDpŝ̽0�I��_���K�L�LB���&gP�|�C�4"e/r�w�a�t*�)��X������-�G��!ls��ُ٤�7���W'�Tm_�����'�W�X��y��];+G`@�cg���PS��%��u;���df�=�g�ǳ ���86|Df�<��j)� �g��F�)�Ks���
����,���ʳ4��Vn��+�L|���_Gf�?�޳�;J���V�z6 �d�HB0y=���$�k��r�;����{f�Jm����n^w^�q,�(��=����������u&����n�eLf�	��c�-J}�/����%G9@�s�z�VIr�m#�s�#@�\JV��}�f�|��L�>��fT�W*�t$���@�o�NK�*+.O:Y�����Z���x�y2D��sl�<�K��s�lɱ�����QY��e�?����+aMF&Z�3k���YZ�~t��z��	t��Z������6ݥ�������r��T���ג�<�ٝs�����C>a�5��X����Pyc���l��"e���ӃαL>���y[Ι�|���l�x����X���x��"�9�2&( $�D1'��N�e|�"ߐ��B&��̔�,Rz���	�N�;��)�eչ�+YIIu{�v��g�~�;������wx�;B����QJ��� ���^V,�XF+s���b�z5��`���T��Ehv���x{{+�q���^�d�8��+U�p��іh@��{0�g� U�oK����W�3??*�j����Gu�7Y;p�JuF�,`��C��Hg��X�mڳ���Q������Z�ڴ,Ц����\��u�# P��l����:��m��gz<���Mk�ִ��6(>�_�v٦������l�W��e;�d��c�O��ޫ>�[���>	>9�����n#����cI���J^�8\�m��^?ۊ�����/��k��=֘�<�=ֱ&���.�1k�#<��~wo-cb��L)#�攭g��@&�� �h�)ִM9g8���s��y�Չv�Si��	��q�{��߱���T򤪣U.��{lKx�!gfB�r궲Ӱ��O9ѥ���,8x���3ɑ��o�=��`��D�^g��E�9����[�A���k�A��S��6G�yϟa͈Y���Y�g�#L�U���_d5���;6?�ʮ�+�� }��˟�����Xm�������1�.���9j�|ͻ�� ������ ����m[�w�y�5�/<�����dj�۳���G~/E�dV辙�G+��Vh��;B��d3 |4�d{��<�~�sc1c����r�/��	��];�;��U��;���J]��<��,d�I�B���(�t���3�%}����l��M�'�`��=� ���}]v�"�"s�:4��>�L4�6k�9f�����YL���ȸF��3���h�j�lP"??��MM�ӏ�ǒ ����@Ǒh�p��L�;�=�{��?)c�Wލu��;=b1Ϭ��w|�^�{���d�D9{�g�$J;�Y�W5(3�1�������b,[6��S{�\k���p��yGd��u)%SL5����1�c_J�6��Qwq(ʎRVs�v@ʙb�ǘ��{M1���H�2��=F�1a��͢�CN*��t5��� ��I��$��k�n���s�����H(��a�5LÏ'�բ�=��\�������� I��
 b�g��M���m�̲�l��D޻R����S�dӤ���i��zt��R���lã�یE|���@�f�%C��O�P�e֮X�f��r�/� Ѫ��m�:��i��^3�!�l`�N��Ā%�]Zu���UF��qKkV{�U��r�j9�7�:�5�g��+��H��ư�I���of�m)����(�{� )������߿��W0�����A����<�|ƃ';�0�i������S�s�Ѝ�M�d: !��BE�<P�\�m��]Lܩ(y�Y�� �
p(u%���9Wbf�6��{�^�܆�1d� "ç�=��3�)�!{*=�۶�7����V[��+K��%p[M,�(��eƓ[�mm��=ez0��
2�y�E�7j�r�	�-l��:����8��6�# 1��}GlȪ���W3!��o�s݇+P����:3.�5�XZ*��P�U�����!�;˲�3G��-���귾_��{���������?��[���Y����gz�ξ�6�9�W w���v���Hj ���p<ff΢�,ڬ�H�;����ÕX9T�/g��8��"�|p��E��:�loc�+��q]g�뀣߃9��� j|F�6��<�}��Z��X���w�-�9�ԯAI�?�ב"�"w`������(�\<��;xB��ϐ/��S'z�xS��0\�Ť��+��[j�S>%�jK�V�I�%����ލYJ��1bw�A���,ŃR��"�bs�iצ�����ep�߭�r��1`8������[E9��}�e��߬����??�	�/gDo\G�z��wҖpddz'�.L�s�Ѭ�ʣr
�@�l��9���Y��ZWdu" p��t����d��3r��:[ζ����z�����y>��xܷ�`~���u�$��ٴ���2�fU�W�w��>O�(����#��f�����r���`E������Z���j9bf}d�+�$������Hf~����s)S��\�����\G���r.�ea7ey9�������uʦPדQ6D���ˎbA:�z`��7���:�x;�Y�u�Ώ�eS+د�mV٫2i�w�3�Q~/�b��� � ��Do���Ǭ~�ڶ����"��t_�b����sn$�`y������}�?C���l�+�X�fG���;ޗ���wm=�%��>+t�a�P?+�Z�fl���bd�ʾ��f��j���n�ɮ9�di�U�#�xh��4�HU���5Ii<���;�<�50gr�͡}>��yfO�~`F3����=�'�Ę�h�u�삁������j�L�ɽ���HV2W���T�;YI����X'�����O�ч�����8�j�|�����򶳞ݚ�Y\�_�SV"�9W6����T�.��f~��x�D�xdyrS��Ί{��IV��8øJ�'�����B@�r��O�7����9�Cn�l�G��l�]+��fe?
����y��H��R�5!����S�#��9>Rj� e�Y_��I+t�\Gď� sd���3��?
O��T����#d�o���9�Y�G�e��p�s{-[��wrUl��ùd�[�<����ח��r�8��A"�T�r�\��^�� |�tdq��v�xe0?�����~'���|"��.?oa#�ݝ�@�~P���=ٌ.T�z#�\����4���VN�V�����b2��c�NNp�8TJ�*[}=���M~f�+Lg!����~EV׏@�68*C/8(1p���%�*�̂��C>�p\Kٮ3̭�c/�h���4g�$K6{�#��p�,���;���9����������ڛ�3����X��-��f�wv�����>��l��pyG�t�u��o����{f�s{ƣR��������?��$'��?����Y,O�.ior���ݪu@��̟y�:��=�;���=vcI@a���w l6̲�6��=YhqkV�X�&������������!�;�(�+ܩ��t�X8_��N����|=Y�h�q�h��Z����A�8hG�Y<3�b'9��9�9���6�A��ȷ���`��30��<��X�8	r3�(z�~ֳ��ؒ�3)rC���l &@ٿ;5��h����٦gɪ��zV`������t晢YG�r�%�������!����y�YL�3���\9�Z�����v�Q�s_�_��Ia Rvum�¿��������y͜���D a�� z?>�q?��l���a��3 ��ݥL4fU�� f� =��F�m�~(�����$��I.&�����_V���9l�!�B~E�s�sbѱ�h2�+];^su`?*V����\���,G�k^0t芣���[����+��ᇅN2ųg��g� ������Nm)�C�У�?�֭䈵zD��k�˗�9s[���?;��w��٭jV�z�N0�fN��w���l��}�b��������|4w� ���(�����&ZR>��x�o6���su����Xؖ�j�w�����r�ǚ�Q;f���j��|p޹����;��%�/ۜ��E�KR&�y(^�!?}���̸{
�� "Ā��r�q�@�z�~R��ų�/B��&wE�NrM�{u���� Z(�X+^L8�oν7��y!�XSp�ګ�͋1}����!sS��,�2"+`q���ʓ��R�6��a�QW}?oT3�pli�kh66z���X"n�[�>��3sA�)��+�G3��~\�P��z���L��mD�x��^�2��z|
���=�L��m[a6x��}4�W���5cV���2�d����^�δA��N���ա_��>�����4����;Pi�߲�l!�X���V߾�{=�������f՜Q�+Vb���nm�w$�Q�D.?��қ`�����*@���p�;�>S�,N&P:��N]0�=��@Y&��Rߥ� 6з�N/�{�x
=�������E�{��6l���V�?�#'�aLyW
���y^������t״2F�}*>�-��Ml��3��ζݺg[�g[�ހ�dN�5�K=0���-`#A����Pǜ�^��؞���|�n�����e�s�e���>�3e�&1cR���쳙�w5>W,�s����{_H�m�٬�e�˶��jj�m�`k�yJ�s����������@[V`G�|�=~������<����)��,Wϧ����9��%�����v {v0<�L��n�+�Y��{~k|�ϵ���UN����>� �:0΂���`��>��^^8�$Ǘ̵�|�<Rl����\�
������@�����k�x�{��u������7����yd ~��q�{���]�^����I�#�Yޑ�& r����s8WR\�q�m[� s�eκ���-�P���=~r��˘L�?�&�������q������6���/9g�k����<�(b�OZ@|o��8���YG��N�%?��.g��v�;�mۺ|��w:ǻ<�h�S��n�\��@��u}{��f,�s+��f,ΰs��ڀ��V{�&lpl�o��+��T� !�\G�&7�+r�$�z�ݦ�fV6� `�ځ�{�}�ض��X;2��϶_����$A��}���}b�X�D�7��G���|S��@Y���pg�̣�5{����k�Q�.u�J�˵V�zW��[�1��k�[u�ֈ�u|o�N�����/+u��jn ��U}�.����~K��sƯ_��9���Ж���z�g�#���&��҄� �̫����}��C��eʥ�
˛��cC�����ȗ2��ꥹb�)np�G���0�.�eB�*=c���;^_�a�M@�j�[w>�L��A��!�k*�TY^%0�Q;o|���p8{��:���7_VY������*TȌѻ�ư����?��j�^�����A���b���0�\$�kǿ5�_�Y���U��{J�H��㴪+phݫ�Gn�\�l�Gg�yf��@Ҭ��u��f�=_��P��/��}i];D}�gm��l�#��9�i]��^_��e�$����y��&��X������:к͚�8^�s�_�Z�������$�{d��r{��9 �G>�On��*�  �;������ _�d`�h����P�TfN/�\��e����i���������vPb�&1 sj`4��ϲ�ge6�,��u9���'���PA���x���{�=W�LlO`J��	��r�ߍ���0���~/��-�ZJ�f��B�6N�6yf �7�3�b�,������~�>���14����G�ov��[�$u��m����9�5��r�l� �!U�!���>��6[��x{{���>����)�@^�X��d�W�ٻ�����e�)���X�K����*�π����P!���´%�l,��1�q�G�FiC?�dZ6�2]�\?�Z<����3��f��c$h���b�:n���ɤCfuz���g)ӣR�2�4�09{��|i/��5���Y�)��A�}.�ʗ�0��CF�:ZA�89��2�th  �p�g�8��ӔYdfR���w@�@�������Ԑc��г����D�=��˫��a�46��Hlr��^b�G��4&��i�HOt))�4�Â9n�Rş̍��e�����nf,��ƺg$�h���Z���8+���&A�YG��#�V}˲�ZfIt\Oi��ipơI�V�<���l�fJ�m	t�8Ѭ��\��zFV��H����a-Gm� �L,����4������q��n>g�W���u���&Up�pC�>8�0�Ծ~��D�yd_l[o�!U�to��U��\k�� ����X�H�L�ll_������m��L=�;�4��Xj��K�2gI@y�{��EmH)R
�}����d�28�1��w��S��� �3�sD;�S�95D�>� ��ΞuQ�7r)V�i�����]�X����,��}c֓�k�D�@)�,�t=f���؜�!GA�-�B���Hן:��|T_��瘔X=����7� o�Z��z��xf�]�Q�*VRf��J�AGn�6]V��ش@�`�,��y�m[e"$ �s�
 c�J��3(��� (�`Q�7;��d����:#�5�9Vp�����V���att�������e�"�.�^�m>h�ː�`#�ݿ�~\����^+a��U�PO慄�������ˏ�s�,�%-��5[C���=<��|��>��#��r�%Kj�;)�����M�L]�m#��)���l�ƚ����É�i�|�|]0��n"53yU���З4���'��<�<�e��rQL ��`��#���r��&�w��;n���S�5_90�O~�Y<c!�zz�qJ{0�A��F�r��	n;�n���Y[	&uR%I&���l��}�٨GDn�+���
�jP�;�8���,��Ф̞�,�e�� m���4�6	,�z �����ڨ	�,���^���������Al�^��+uj��������@�f�I3�N.KL���
����R�%�O���l�����9ǒ�$hK�&$�t�-�}��&���� ����2l)&�b�N|լN��(�
���+n(�����+n������J�¢&�]N�}���h�s�Q޹�)��~�|�Mf.YqXU�S���@/-˸F�E��(�B�2�bxjR^����f9��^� @c3O.h�f~�)��m�V���,�z��w��N9Zk�H'=��#�\�9t��Y��>sY�:�A]�C]HH�ӇǙپ�)[~f����b3�gK���音2fm��,Vl��{��b$V��Y[��X����-��T=�-@���D��h�)˵y4�s�����hǝ�?3�c=��g��,@rL� S2���=���pc%0"Vzd��z�e�g۶��#m/�	�kB�Ms3[/����dNu�iҵ���ȕ�S����gh�����D|ٷ��S��2o9_��N���n}�v{��=�7'�A��$pI������{M��O&�$#����s����A�B�k��2RQل�\���q�*�'=g��<<�k*�p����
���O�=Fl!PX#(`|�.ȵ�9+ɏ��m����+J�ZG�8��ԧ<��ii���y��v(cV�v��r���:��|��Z��:(>�x�'�|[7�LYE���1�9�v����[}�3��.C2�m�o�g ̬~+N�F%S��t�{����M�m�B���?�#���Y�e=��������jC.րnU�l)��љmV�5�fm�y�>X�Y�u�{�,Oy�hN;z��?���k�<XΞA�+��zvB.��d�ˣCQ뛶��g��{�e�a|�~�k�*N3��f��M��k�@�L��<�i�����;���9��_����淂Kl��H��-4�PO���7�ܛ������������ƈ\�̒C=��&u���>��|]Ɵ��R��0ف�gn��C
��\m ����7L�M��UQU+D9�j]?���5(������6�C-_:>���>�sL�EW��b����&+��9�CP��XP����6�c/l�^���v���4���~s^���hpq��ifP�K.�ᶵpRv]Ǖ=NّFo.�y%;�ݾ�4���dX1p��}�|뚣Ì��}ֻ�1oW���Y�<��!�2Z=�޾|�%�>�>�֩v{�#�X�^�\��}{�5-|�;r��f �Z2�+[ɜ��C�Z�=7�-����!�h����ƃ��L�>WO�R���ƶ�\�ԃ@.�u��0�Q�ޒ}v�1�?l�	V����� SHΌ��/Kr�1rV�\YM Ⱦ�!����R�i���̔x�,6)%�n�(�����O䜱scQFCk�l�n����.��������b��;_M�pa�R���/v#��`�@��r$s�z�035��|X���ɌQ�1-���Hj�fVבh��Z��a�+L(�Q�J�X^�=�f鲸���Z�Q��Y?/]�����hmh��V$���Y��\2NqϪ�z�b��mׇV�_,�����78&�Ӿ�{{�(3����5ZV!7|���_�!|`V����iJ,���� {"��F�.S�e,�s�[a2��\Ñ~�%�K@�?���k/���$�
��!�`0sE���\��H*��L���	.�	�v/3+�;n[�
o����i#Z���X���Zx�8d��� ��sK��3��ƛb��l�2�.�^���~昜}7^�B�*�f���6Nj���{�I�ƙ̥���ܾY�+��R�W�~��^3Cr�ʰZ̬t:���3�E,$K<;,JF������b���qV'�[{G��.�/��8��6[��pR�q���}��e+�ҰF�m�Ҟ�\K�f뾎k<�H��U� �.W��נW����>�(�cU��8�p�*h�Cbiېz琽�@��L��[)\T�+�ѩ�Ĉ���ߠ��LTv���_c������K�Ql<�d�js '젌�S��ݯ�u�'#挈�qɴ�{nc��4��N�Z�B�vuCՋ'�D��q���е]�c�	��+9���i�G�8��]%"��gY���vD��f�)?�Hp]��,p;�d� �3��MI�p�Rm5�Sg ��{�T��[1QmlgHp}�]+`������긥��~�{=>��_�5S�[���V�]�Z�f�c��eh�~����@?�<�Y |��1*���H�嚕��x^��FH�Y[�K�N�	 ���]~��Z���¸�����#S��Xk���i�R�L�a�:��2���h?���{�v~�m�jb�S�}����"�:"�8^wݗs��F�c�KPv�Q����ɣ��1��B�d����K�d&J��3;Wq���+��4��yWyL0ç��h�b�"|r��N߶M���fʿ���B5k�#�T��H���QP��K���>���\�Z�y�B�W��cՑ��^�9��U�FC�D�F���	ĸ�uM�(t(��8;���k��j��;Xgh�2n�۲�G5
�fie�9��C���G�,�͊��=�]m���u$����>����-�ri 7sHl�6��U���gz��YN�׶���ڔ��'	��Y�,��̽ֆ�����J�u�k��Sz|8�C�z}��암��2Ey���Ȍ?-�y&@�3`/�����_�]N�klL���Y�y�`���,Tu����m9b�A�������B��a/���;-+�y������n���ZY-�þ���Ǉ�#�C��ZtP��8��X�dN�wG�p%<��H �+��*k�g�G�<(��t��M�#E�`~t}�4"��#T��%��Oytx�>������l\1�imU�39z�� 1��m%� b n�$&���,Y�;[�q�d��򯊶K<:X\a���h�l��%c*���4��#��f���v�l�	2�d�]7�%_�.ψ{BB�"1�A �����u03�_k���'E
A�rΉ,lT�:>�h�'��޳���ZF��<t�W�^��I[��`�~�C��S猪�3�mq���2�ޗ3&��Ӷ�[J��$�Շ-X�������ڌ�;�3��f���g�G�&}�T	���m���>��_��6��X�T�W`x&W��f2g,,��*a�.	�Lz����j���0'���7�)�{{\���朼V��7g�Ԟ�"m�mь�L������Y���/�3z|Y̵���q�>��^�/��9�.���L�;����u�Υ]r�0��F2'��\΀s-y�7�/�	��@�| pY�"hQ('� �G �c]qr�8�P�CGA5�����Gv�Ԃr����������𡜾���O����� �>�D�������q��C�_�zMz��OU�Ǡ���Z�8?xZ�K���~�������
 ��&�J��E2�V�dK��Ǭ��d�����y��nMe/�Lf`W�ɋ�;�3	f�a9I@5۰W���d���G3�d� � �Uve��#wVf��g���C��@�*[n����	!�A���M�.��c�ǰ��a☩���@����˺t&�Yy ��^��Z R�_T��<�5y?lD
9�='��	Ⱥm\�|��zs3�S!>٫�h�M�=�qԟ��3��^�T��u^�;�vz�-��;�������)&��������9({����SQdcˤ�Gʎ�H��WL
K���nc��
'�"�	���<�
�B�h�*��^��%ۡ����.S�C�h$������y���Z� �� �Q�ҳdH�����o��wa3��A�be����Lc(�k~�6�jU��6�]Þ����m[�������Ҝ�??	�gzc��:�&�����+������ ����H���c�u�W`�L�Z[ڜs�XD٪Ϋ� ��۰m�k7����s}�vYF�=��{�K�D�}dS���r��e��>��u��u�v�����TD��k��n�CL�o6���_�@a�xv��r ��S��s�P���8�wvȡX�@�Y���չ��@r����%�f��3�O�)���K��d�����P�s��Jx��{O�s������j�L���aSt)���=�>C��<�E4�\���=��1Yl��G��&��r6��;�]�/��+[N	HR���s6u+5��s�iIʑ�V�AmL��+m�be����Gǳd���K�CjYrtP��ɢ��:�?�V���w�|f�b�uE��DNό�+�Rkc���Y�M��B�#�	'W߳��:��ƴ �ԷG |͠[*�S�[��W�[��RC���}�u\q:P��a�ɪ���3���gߜ��e~m0v�L 
`�ۆ����#1g8����)r{��v�!�����an�[�� �`�$ȜQ��;���+U'���(�ܭ2�e�S?�A����	�����S�J��-�=�x%x}�iG�������PJ<����3[a�x!]ej�R�Z���������M����g��f�7-gA`+�ز3�F`�=R��0J/���f6� �d��� ��w-}k�G̦l������@+6S�����#�߫9{u�<��i�����6zV�9=fR�}��<�����L-G��sm�k�V�m1��a�{�|o�Ѷ�O}㐑�:�RU�{��	����s�|��#�ui%�gn� b=Bض[u�a&��X�d�q-��\��;b�#����v��N���x	���&�!	�7Ǌ�M�\p,�����Nd(��h���#�O�L�]c��g^��
1�!#���Wm�6�Ҏ��y���-�s��i�+հ����L��Ih3��R�_���N�#�k�����wFM��CM���8���C���s*YRK5�Az�z���Vز�DA�syhj妲��A�x�C��m�m�[��ol`�qvu�@�����Zu,�:2]���?~� ������`�Vl������8p� ��<��7B�of���R��������puW��^w�3�D3\?ќ��g�R�l�9�&d>*�8H��z�m�w�SN+;-l��3#[�J��!��WB������B�2sd��>u9@�PA�A�' =Z�%E
�6������Bj85�� ߌΟm�+�&�5g��S�U�&qV��4��8�̼��-܆f����A����c�:X��%����b0��3=IWL�~�Z�H�W��}Πr�<�vm��x!<�ls:�y0�4��Ȟ	=Ň&ma1��69����ׯ��)d�K�&s}H�A��gz�u_k��3������Ư�h$�[�2��㰩Sω���\;������)Sjp�]���Y,���<�d���a��&q9εز�kf�z��(�m�9���tl&��s��/��<�9�6��q�L�B&�����S���FU��s&���c�Y��{�)����m�N0Z􀞩��ʐ��H�"�Ug�Qy�v>C�Ƿ�z�\)��`�6^8h����G욎���7�m��Sx��d�Z|NtY=Vϱ��;��=�{��,�_v����/���Ȇ���ش�"��t�&]�l��*5l�w6;�Z@�ꆿ�U?<�5�be�i`�iGZ��6�s��#Ś;�Fr� [S�����G���{&� ��Ι}��6H`��.��$ᶢ�=���wpF�"<��,V��rЬ,<t�8�S��3�M'eMJ�t�ZX��L�!l-�h��a��r�����3��u�H���$z8ń�"¤�X%@`wTʓ�5��Æ�2c2�.ң�`4g��:c^�L��g㉴-��R�m���-�q6e���s��\O�"=]�u����!�E:��
H�쏔"n��C�|�
�7�U��)'F*Lc�]�|�_VY�^�/�V�m^��- �b-f����ɚ�R�
 ֐�Py���v�2��,�<{��ʹ��[2ca{F���C��\�ݣ�e�Q�]��M�\Wkޕ�֚���g��ոҦJzav[�����Ɍ�9K�*׍3��L>Pf�P�� G���+�z�2�,�D���wp��{����^^��pǒ�\���R��g������)QNde �"gp����jO��&��璲����+Y�qgU����b<�Nh|�k�Z|g��Tf횷e�^�������l�]=oˈ���m�������"�c��B�e����d;zv�d�r1�u[��θ+@'5�rs�9�
�_��Y fƎ���x���9�J:	�,0����g��Z�7�8�g\�M9�΀V-3�|�<Z�,������ѹ����c�[ ]��g��=�k g���H�������A����Dץ��,�9�����]&]GLھ�#�͋<��IH����*S��;p
�� �iO��9�@I��_>��8�E�h���(�N��Q�D�=�o�9Q;#HZZ�C|�����=��\vp9�������;b��S��~/�Ǘ���1F�n�:V`3�\������A��D���:WJ�����_!_'%W(|;E�b�����o�~�;�}'����S����z2 �Y����h��/ۭ�_/^���6]v��b�1��y�z�)p\(��+�T:-p�H�8��<Ru]���ȶmũ&c���l3`FC:"ͮ;#�!U�Ɖwٹ��\c�g d��ȍX�uVG�)Z>2���!�Xf@T�����b6��m gcwV?;�XeKF��XG98�sʹ�/W���?3���X,��!��X?���3�}䊑�u�9J3 ��΍v���Ɋ��]���3صYh$�o���(��S�����{��4��m��~����Lf�֗%P�+ ^�G90: �ڊ�.�w�/�4Pb^R^���C���K��N�,y�!�>$�i���yme����<B��U���x}}�O)UOw����"e!}ԟ���;���z�]ԟ]���g���\}�,a[,�t��Ң��{65 ~|1� ק�|D��<������
�?��"�0�=�?��j�Df�����q~�9*Ue+����}�{��x�5<�C7���x�T�������@�#?�{��<q��U�]�DZ�g�a�a�h��a�D��~?{uF����؏�������n�4) ��"yz�uR�-T[��r<���m��&缰��&%��u#Q
�Lu22|��vc��i�|�L��22�!P�)4�V\�Í�Z�	a��K�I����e��2����@Ie�ᕊ��1���!Kι�+:�,y^�1]]���g֞U��:�
�v�*�Y�S��Sj!.��W�v�hq����A�$�?��0�\�=$H�?�zH1�g�/�Jf����M�S�R�ׯ_a���WZy�b	>�5��s�qm廚��Y�9 X���9��wZ��Ȳ�<j�� ̜�,M��oN�*>1�,�̳��3I���r?��8#�H��8I`ƸS��,��]�\����^T�ь�{��W�o�����2~�^(|��s.��h~�Mf�˔��#����>l���b��]  Z��f�'ǟӭ�yMN4�3f!X�#pk'��������!"#�f�����pR�@z}} Ē��W?,���R�\9�j#}�Ŧ��2�>�������u��ٴڛ�3��6��:��ղ���沼h�u�C�s�^����b��v~��rؓ!m��f$��Ά��S��u��:���g�v� �#@t��?�S�2X�� B��V����%Kuj�m�7^�_yp�����Y�g6���6ڈ�2�l�-iB��C��r��5hvm{����Ag�׶��]��9��"	ӫ�N��0�o�>��`��l�G�NmқF4��{�Q�T��m�LM�#b���s���X¶�N9�s�K<w�����ة���r�Mw���0�!a��׍���j�A���gF����g�$�~�|]�4�:�0�t-yv�2@�i���#W���v�S'O��5C�O6�>x�gȬ\���=ֵ�/�������k�?�];��g3O�H��:�DZοJ�s��<�}?g��MDz�M,>���p����������W���lx������~'{�<�27z��^�� ''�k�GL�*?"������>�?ڦ3Z�����|Z�	��� ���3�u�jn?{��L6�Z��l�M9�j�d���̂���%�@�Z��=P���=3��,�N��d�;�|K������,U�ݬQ*.T���&$��1K���%_�9#�a�>P�HRY{�L/0��|x��y���C��w�! b��b��]ur H��L9�g*��-g�q|�mDg�}����k>�^�Ws�T�m�&�`=�����*��Pim��<g&���|q\�1ʶg��䵂{�<2���:m��F�`ł�j�m�6;J �c�ڢJ9JO�Ǖe}H��zr-����#���3���(��r�fީ}v60���~��9,�)�1�I�wd�V"�m9ׂ�K`6[K���� P��X{ҕ>b��9��3�w:d���D������[�>�9> l	����=`*E���^ ef�R�,�����0t�Q����2��;1�m�f�����%��/2=�#��T=�k�ɜ�5+a�5�a��>�Ӫ��13}D�f]O�Q}b��-��._�,P9k��Ŕ�� P)�v��s�ƽk׌�u�NN�x�]�ӬQ#�����m�UՂ����[�$��m$�	�1}�ʹ��%x��0�4	H�w;�������{zvfC���?���R��Bgw}������g5;E��R4��p���rm3�3�3~3B� ��l���YďL�;}
��_iAw8����ؖ�9|�~.k�\[���r]���;|�u���Wei�ZE���BVI�v����\罄,�1��N��d/~� �Gi":`&
ɔK�� 2Kˌ���)_d��&�s��v�
w���ȕ�,p�.2���2���)`.�H��Q�J�,z�tޘ�Q�P8��,�����	���+�1(-p�R9�Ĳ���5�:��cU�X���ޫ?V w�vg�믿 �PB}�v�
H���'�����j��y��:�NlU��7�Y�VVB�抚ߕM�P卋���޻�ns&R����b_���-�*�K;����W^۶J��[�}�]���Ǐ�x|}}��0b�&�A*���G3���m�[:���N�ȫ[���㛲�|}��@��������62�9ܭ�%����h�י���>^��w���W���3����`�����3L$���p�b<�����-��kc��T����C�p��k7{�kpɌᶅZw�qG�(��E ��շ-������)E����<��f�$2AU�@�yt@i�i=w�"|Ƹ��A��&� p١����lO/(�H�_��fg�_���Zl�;���&d2���Dl�'������@�Ӿ!�O�_I��}Ev`g��UY���-�_mQ�6|�^K���5���Fut�3ߗ���i}&@3���F��:S�X��f��q�%�l��l?��{F,'9'u�����s�W�hk�>�y<k��ƗL���S���X�}�Ac�6�BتɌn��e����u�-�������xNh09�+�=ͬ�n�YY���K U��h��N�; �%��i�Q�=�q����~G��e�y�l<bm)3� �#RNx��v�~7��鴲�Ќ���jlL��mCJ7�[B�	�m/�k�ʾxGt�Bl����kk�Ėɾ���3X�J5���i�n�����Q{X����3�a1�2k	���m��y��{��g�3C)���j�E��?j�������I�g9i��ϸ�G�7����^��lπ�h=��{�A|v�JPc-�Z�Ξ�lLH9����J\+۠�j��L<��.�kʜٟk�ȑW��?�ЪY������a�l��s%?��:+ �Fk��� �\׬�T���h'x>Ƹ�~�#&Y��S�E�dZkkۼ�Ke�A��$�;ʗ1���ךĬF/���&���~�������'ft���:�ɹ��������z�Ґj^	4�gV��G���G^3��Ұ 1]��:�>��𨍭����e+������a=���2�S�6HG���4��*Zj�\ g��ʶs�ʻ"h6�)����JŁ�Y��_�^=�
t�<��=�Σwf�oxJqe��K��,��R��?g�=�G��߯+��s�.y�՚7��._��G�5�=C�=���KY��ה�3�.w�V��T�m��7nS�	�]�z✫�y-�=�=E��!��/龶|'�"�)�e1�ؙA�Δۜ̀	D�=���c�_HLk�u*�
.��H���O^��<�  e�ML.޻�M�ۚI �q�h�u�m�=�T�L�4�<�A�q��}g
	�t�p��*�����Q+P���������rfz!�X|�Ŭ�<;��\=zo����vY2�_���#���􌴨 v�"�α�M�q���%�:�������$�����1-ݕ��g�d�e�6��6�,��'�'��`�'{"ρ�W:��w�����$�Z� �ϖ�1�l��T}�u�x0���-��;��s��e�{����?���h_��Q}E՜ ��(q�~�e�m�4�������?~P��\>/Z����ƀ尵�f�Z���	 t�~?��e!�H:^���������ؽ�3�/NA���U9^F�O	=�������Ŕ�P)��}&'�jBX�C	u}W�ha�m�zs���N)�`�q�>�i��&�k�_[y��<]��;:�H0�y�^g6�g���H��@�m�x�&QJ�^��3j����P:�u�U>3��!�K��3c%�{�7����C�i�g����$g*����x�!�ք��s��/,���1'Rw��G	6{��Vw�BO���g��<�}�w6��d*���D�Ô�R��9LٓҒ�=ʵ|�q�e��(e#e�a�B����՘S ��cY��we��)�N��N�}W���{����=���s�bbU�#A2��ʬR��J����d.��g��u]-�FoC��V�jZ����6i��c�{>":n�Lƅqf�s�Q�lu�Up5K��BT���t������\u�ь*?}��.<	��l��Q2�Y8%��=�{Ӓ����,�d9���O���t�k�����Ϸ��d��,��8}n���� +���~��	0u=2.��n�{N	ZM�fr%G�|�6�2�{�3EޫR�4.����>��J]�U������L�83�I6�:��w�/����s(ES��̆��XD��-��M�{ :�&���f:ðг��#���Ł=�6�d�MP�{o��j��s�]��bg2�ݚ�X%@�m�"ۤ޽��s��,�a
4P� �Y�g2��ܨ�V�V���}��TzƳ���i��>�����J���3{T/����wh�W�<Tx��k&�J/3s��G�s>86�t�#�;(4YS�����̸m�<�l%r�����Ǫ��9�:�-g�\�nXk%����	4�>��T�[뇱�_���J{�#q�e�ε�{
�N�X�]_������(IT�G��Z�K:��q���% ӱ��wH���-p�e �p"�Rq�GBH�>;�= ����)P�#������G���sp�#�o�����k���y��q����gZPSL�5�U>�ro�[��e{N�x�<1�	P�v� �ɀ��7a��X'����ǪSn<��xd)����s����q��YE�t�O�#�loDg.Yﱺ��V�Ij�0��(�P3�|�A�V�o��F�
�ȦԺ_:itkc����$[x(h6Q����%}�j�f+��m�?g�晪b��y�m���fdǔ���vI{������ϊ~V�/����;7�Q�x��!�w�@m�_k�����,>�|gE�Y��{����6�ٲ"�\m���j��y�; !��_�鴣��t}^�r�P�35S��4�~�!�$ (�$' ��O��99�OGN�Z��~����=�9;�x��@���N~�27k�E����J�z��F�/���Z��$wdd:����a�%��(�hr�d6��&~1�r�6e�`���9�h�o��4���S"������hm���E[��Z��K��]���g`k\��ޑQ��3����6I���d]3�6�0�,W۠C�h����υ��B����&	�w�r������rՀe2�w�J��#�,�G�΁�M����{Z���̤�mkA� �#�D>9��4'9ۮv��}y��z|��Z�7P�!���i�͢��Gjs��)+��������-��s?y}�{��y�Ҿ�^h}�@��"���;Bx}J��)_��H�,.[�e�-��l���̧w�|"����X*��״���kU� x)'��D����*�9���۠[Y�nޏa`,U�%G�Mf'z.d2?_Vu�6Y�YP6��Ȱ=�e�Ɯ���fr��,����G���,c��١E��%���8���{Vy�M?��UHK>T��#+l3�cȞ��)�h~��6� �3e��J*6�M��\o.q�,���9��;�q{F���Y����=ܮ�����[ڱ�ګ��~&����΢oH�����y�Q\�\nOnW��\�Z낁���6�rp�E\26�0@z��1ה�,�I�Gʩf��5>Sa�DQ��o<��#ȳ&sc��~�<]���Z\����`��X��g,�:���l�l��Aě� W0�X��z���u�L}8�����Ԓ�|�]�x@�l��3l������l�^���ۙ���#I���,0y�~�g�v�������U/ϡf2�l�S����m�##��s�:���8bx�6����m�u�f2��tŢj >@����,�2����9� �wl5WR�$R%�r�5"OJ�����w����% ������_�sp���Advp`%�w�~�ȹ0��� ��Jݹ���9ռ���#���z2�=�����������^��~}}�m�a��٥��0���a���=��M��d�lf�5��!�����z�zz֮�r���s;�{���<6x��S�L$ ���@�7t	�x�36����Ϯ�s�31Ɩ��Ё��G��Jϴ�v�v[�<��s_����<�>Q��t��޴H��L_j��
@�����^��M-��tCW�V{�22����>_�#��˘��s���+�//Ծ��ޕ���Z��4;h��Z;���?�OG[�ۢ���_kbP���2�ӯ��5���o��>0��<��/�d.S�\���m�W!����J/�����}Q��l������vk��,�ۑie&��}�(���5G�% �?�������a����p���AQB���3�w���s: Vμ6�����X �0)&�l4W��g� fu6�1���Y�, �m��bt�Yы���۲-_%V�b�<X2c�ya��-��a�硓��׫��<���7�4�r�%{��ћ��x4��ڎB�m0��ka���6kƽn�'3�<����K�q�U?�q>����,�aX��䟳�^Gr�\�rΦ���v|��i�#�]��xM������#�%GDȘ �Ş��u������}����𘲶N�=�- �PcrgB����A&6���_'h}]��O�Y%ǌ������ 2�#;�Y4�s�paC��߁(��N�=>��0�	9&ĸù�=��-����\84��I��2����<�Q���\���5YW�f�^k����ڳ�^�ᙛ�w��������|p;�cF_/��\aѨ��V�Y����G<ع�E3g �W�N3/�~\�K�Vz�sV���#�H(�𜹼"G6����h����sBp��c�c��Z�V��� �m���&�-̐f��_�����m������� �~�����r�ߛ�$���="��}ϸ�n���-R	�����ZJ�3��r[T0'���R���% ����?��u��ÿ����_���?p���=���;��6���=(�g L
e:!�3�`+hgb_�S&��=��X�Sؒ�lZ�%�vb�����:�|6V��re��,>�����ӳ}|�>f���Ϻ�b�f�|eS�1���wg@��-2X:�_b��@s��H��AZ��a}bL��l�7q'�V� f)v��}0���r�L���?�g��s�Ѯ58}�����Q���?jw+c�4h�2n��Q�usR�uO�!ql�����W�[��=�!2���z)~��kvO;�Z�j�T@ �xr�	Td|�ϐ#�w��T��Ƕ���q1�K�I\�=3ʔ)���S���% ��������������z������?�?{��a8������g� 8���@��P�w�<��K�t�"!���u��m��`N9U���ۆ����9!"!��#�Kp��k�?~� @jⷷ7�n/��bL��b\�I,��5|?��0*|?��&�ft[n��!�͙����T�����K�=kÙE��:s�h}?z�[��I����g�Z�po��;��};>�jSo��13���չ�.�n*uV���^�h~>�����i��m	ge�6�X����g�~�ƃ=���X;�H2��>�-�3�w���+�/6�<�)���)�a�Ƶh�Z��z��;Cz�FAjVx�.~��cUg?���k��,���<�>�#�~��Xk���+����V�,��Z�o���w����D�l¦ɤ+�sy]b��wJuw��;���;��B��ϟ��}/{�{�����,�^__�r{��m> �#;���9xW��>f����w���.w���g���������gy��|{����wOO1���tn�\�ޕ��	>��G��	
�
�$Y7����Ug�^���g�䱘Ќ�m�޼N��Q���
����L�����~_����U�___b�Ny��W>��J{�:� ՙ�q��1���h��A��Y9�w;��	�6��s�އ��Sw���l�b��R�k�E}_��U��g`�
\>��!�D��t5@=_K��g��l��u�]��H~.m�%c|PY�ź_~~#Ӫc} �9���3�ϒ3��s��~.k��90;H�x�%�m6f9��}��os�c��c�+��'����C�!��-l�B�?�ߑ��Ӷ� N�"�����V�a=�����]/��A�G�ފs3��@u+��w�/�o������'�������_y����w�e��85G�IL��  |�7İ�L���x�����J�D����wx�m:iΜ���$iQ�d���E�/�=��*R��|�ʤ��TGq�T�H�	 ��ީܯ:���M�# �Jϸ�,�\����%�2��x�^u��94H�՞S@�Fs�8K���ޮr������� Ԛ����5�|U�������������:������{�L��W��3�U#{��{�����B�a֮�{�å���(�of��a�|����yA���ʹ��y�*�<"@xM�!#$_U�g�����Y�N|�Ԕ�Ц����c��gȗ�����ۿ���?��������?��ן?�p�{���>��P����@���6��a21��,_�irv$ "�L�`�V�������Ǿ�u�Nk#e����U��;��Z/�zA�i.��Ѫ[��U����~+l�j�h5��{�&����g�Y��,{!���n�	j��{�^��=fX����cľ�����mï_M��3%~03��s�]}y-|���@�:_�ZM��v���X��{�zF3��r$k��9����c������#�C@��,(&��k�h�����v��ի}���CY&�֞���{�����Nk���{�y�Ǆ
�7�~N'yF��4�Υ�V5u�#^^^p��1a������a3|2�1��S�C��FJuK9�c3���� ����/�����O����������)��*� �p���� �a����0���);ĝlc�H1�a$	��fOAu3�h�$�onP�{�u��^Ĳ�ͨ��"������/^:xߟ$��W�/bg�6lnC$7HY����8�]Rچ���l�&���lum,.7�I8�G�+7��6��bW���;]�����s��f -�p�?gv��
�s�3�`��S�n=�5��c�9��2�}�YB�-�Y-{�f)�Ŭ?�n>��Z��)�����辖:�_cd;$�(ן�a�?���5�����<�y���(�}t����ײ�Y�Ug�������\96����>���VL������`�5����=|��坘�㜋l��\�;j3Am�|q����� �������3�T�N7b��ǔsݦ�����Et�0�̀�1������������/ο;�����?�]U��@6@1��xL�X��S|g � �0�b� E\�z�mN�J��
����@e�����8���,�W�@�I7U�<�F����N�,۶��Z�l�9��3>�hÞ�u��%�v��Qo�;���WA�j�M%Jmm[{{5��g<Ԑ�?�s��Kݬ�t~�KY�kC�m���fq(W����2g����s���w2\���:D^aǤ������s�K��z�j�8k���V�f��}6�V���0�ev8o߭��Q��yo]ۿ�f#;�z<e����t�u� ��DF*�u�F�>o�v�!��r���F\��Å	H�#9�챘~�g�)��~'��(�q���M�0ҒsIs�(�e�=��nq�a����A���K@f�6D8�p��n���v�!�l��6ʴs�m7� ��㍀�N���8�W �s Of8V���$�@��T{�j��Cq�9K�7�B�I��<j;K	F�6g
}�H���h�9s��>?� �ڠ���]_�O�g�Z���h��(ȝy�JB�e���3ʍP���~4�$��-�}��i mIg����92��Dǡ쟯g3�u���V�{�i�UX�u�du}�g�t8,�Gɫ"�i��h����1W%|�=�k��د�`�lN"���O\���Yk�j�~�}���{x��$��I���	u?<�F�P��ǽ��X�I䜋�y,?	Sp����2r������[f�.qc)v�C�}��y�6������� /��^jJ�ߊ�/��!(G-R�v͹1|�])��ː��i0�v�Rhci^�����ږ�>�*��~��e���l�,��ƶ�O청�O/n:��C�˴�k-.��L�� f�Q��wr�)���g�O�ל0f@��({��3m��2�]��~� V(��ٵ�8f�t��>�q^��~�>.O���
�+��Jmf�T4���9?�������`�+���v��v��.�������H������2��g�:k��/�+F�"�2ن���y����_7�q��L���Yh^亽�1D��^��9�2��ɍq��������8O�����2��ڑ>��.�(����>�_-_2���<n ^bB�g���������6rp�e$d8 x�D��6��!�� �y�x~ٜ(�#�-9]N���G�*-���3���k�hy�t�j���vá�S晐"�V��2��ӕ���������T������Ƥؕt��\�e������H�^$q����!8��z��t?}��&��>��b���)&�n�-��~]�L4�2c�tY|�dYV�������n+L���Ϥ}��u�sv�V?[`H�}��ϐ�4ғ]����嵲t�T���֘f��tLS��:��GS��MV�ѷ�r �Y���A=:��$iS;�C�#�K���c��z�f�t��{Ϫ�uڟ�P_z~��к�m�l�E�����_�Q�G�G}�ߣ��
�{����yW��n�.���xف����������!�g��fy/B�pJ� �n羠?c���i<��׿QLl�n�L�\��^��\ƶ9䘰�;���ضM�#v n���G)K�-��8c�2�!�\��$H�O�I�n�n�����: �6�SND�͖�$ ��d�Z,![}�S�9����le�<�,0*���[�u�P��&M[��)�?is���<�9�"�'h��s�Ms��\�{\]���c�ھ<�wY��I=�¬؏�2cl��R4(�11gd�ϴS^sx��g֎��ِ����jd3vg�O3pYչvG����#L�j�>Z�d	?c��T�]�������g���G�~�}�u�������U�s]�!��ŀZ��l�w�e� {	�����gm�y�e/ ��֩�Oi�"����0*�ёX��i�sۆ�vlaC�6��!��g��}�.AdRh��3:����2�:Q �?����V�G��%����p�	�9!��3���~��7x�����Ia`���|����`2A�/*��#�f�֎?��V�K+��>�d!�V����jm�9#2 ^�@L�~�^-P99󻎽��.<�~�� �^D�����k���Z��ja���Θ}��i���<S����Qy6�x`1(l�[��`X3c����g��!���w���!�������n��o67���vu�@�,��A��׋�éTO��L�P��l>��3�D�d }�,�Gyh��������bMOڭ�)Z0�i��?�z^�w�������pU��;K}[���+�,{%�L����n~?�W�̰Q �jgJ�q	�s�wH�%t�̺ö�tze@�'9��N�C���KU�Y��-�@.u\�����H5]��*�[�p�f�z�<}�R��NE��
�����Y�dJ-�y$�Er�.̾[-�36Eާ7����ql7��(әr��w��y����}��E^r���Җ��z����y�^e�U�G�[,�*k���"�����ٕ�5Hw���0�õ��jm������!kV�������x�ዴ���Tȃ����c��u�!���$��l8I�y�S�LV���V�S�7��:[~o���j�p���vO))К� ��i�IRY���q�M������m2�8�9wAK|�D�@�������S�	s��Qs����a#�w	�x�h ��Y�{��ᒃ��*S�@EY����u�Ȳj�E���'�������t��2�:;�ve��z�f`����p4ɏX?]������Y5�<ڠ���#�8K���a�x�zT,&�hc�
j�>��e٫qc�W�5���X��߯�t����,�?ϫ��z�G����e�~���;ڠZu[����;]��=IV�j��F��Hc9^_�[�V�S�_ڟ�uʚ;��T�N|��&��JBɴs�ء66�ig�֬B��@	��*��sF	 ��;��Γ3���_�~�w�ˡ�D�Ƚ���2�I�;_}��dg#$b5��rr��3_)_2�=!�	���"R��<�ı3��ޑ-�󮳉��(?��t�{[<��߶��?a���IX�K�R�����f�O���l��k�~��!�E�\�K��4�LϞ*k�"��u��ʼ���ʲ���\���vh��gm�����<�ժ=m�g
��[f-���~�3���NJ��^ɶ�Y��Q��,��tvZ-K&M���~��5��:����v3P!��1-�Qߝ9��r���굃M�,��5����u٤�|��޷g�̙����t���7�fu���<��|�w	bV�otة� q�#S���̿dZ�!O��:��Lz�yH5_y����i�U7{ ��`3؅Ro�?ﮫx��h z����Y�C��p-RD��:TJ;�ZFٍv��I��L?xVx2��CLi�@�f��: �MM?�^0c�u\�ޕT��Rĭ����g&�n���g���.��t��@뿫}��Ί9��0V�<*��#1{G��|��U{�˘�}�n��b9
��JV�����Z?[?��̳�SN��@�P��匜���0Y�{����������O�������d�������˹���;(}����k@fh`2�͌{�RY�����<A�<�Έv��H��-;�3Aܹ<����}9�v�<��m�����2ۇ��d eY\o�|m)�y��S���2�v������ҘSN���<�M�NX��ؒ���HYlg��׮Sdj&ÐhF�#�ج���j����5��3��
��6�U���{Vu�ur��9�h�t�w�Փ�X1�+��:�1��Z�������K�^]/ (��\��yߖ�
�r��ܷ�ۏ�N^�}�]�k�.�l�`>�蔿�=���}gj�����Υ�1'g1G��|�1S�s�m��o��ײY?ԓ86��iV�w�׀L�|���b{�Q"3o+�	�����X�z�L�,_�P�C[.�)'�{)D��D�S�7S%������6��)L�e�rh�y��,���K;r<n��s��n��j�|������	 x}}�v��T�y���X�j�/BD�E�T��	����Z|+�Z&�d+��Ó]����j�E�aݿ�,l��7pٖg��_#��mC��� ���!G2;@�r�����k�^�b-0���L6�~;n�5Ng�6�����������Ҳ:X�8s��,�������^���H�+˶ �k���g0����}�Ͷ�}>-#Ցĺ����3T {���s���|�v ���S�ȶȝi���U��_Ga���w
%�m�)���)��oW�Y��n����?ѯC9'����61a�}�16}������@&���J�b:f���B�d�)�=��YR9���<x��ڠ��>�AU�#�v'���i�^{m�3]�:9��ԅm��v�d]b��9���o	v�&���T<����m�̹�����L.���6q�	(���0RN��P(r#��:���Y<�:?#����; �ٶ��G�[=��pt���u+�sT�s^d.i��j�.�7.��D����+繻�!+�l���?f��F,�gg힕ԾU9g��u?[(��,���(������N�J)79�������)�Dփʹ�:L�2��j���&���ׄ�4ͳgi��)��~��L2;{�aZ��4��s>(��x���3��0����(�rp{
-�f����/��l)!潂����~�X�:f�V����΍DW�m(�q�9�ϵHݾ�J[L�r�E���|����CNJv4����H�ltuB�q��4d�=�N�5��o�9�)2#��v��b�c�Kf��w�բy溯������<<�i���(��d�x��%�h���� �YM�����)�r��Θճ���G?:.����z�6"�́�Q	4%�d�z�~-� �l��A����BA��"��/4����y�ZT�c��[��q��ĝ2����xo���^�m��Ї�T���r{A��O?G�P
���fR�;sA�N@��1�(�Q�@l�g#�?S�`|d������@9Uռ�0�=ٵ��>UeG�!��:�b�Vۜbw�V�b�͋B'�x�
P	 q/��A ۜ3rd���H�q���ZԌ�X�0��l,��pr�CN�G6ݣ��y}�XL�W�f����{(!�>�fz�L��_��l������#O@޳�ؚ+}���Sm�l��՟��tp��	�L�~4��=��s%��)z��r����-��-=�����5���P�e���}�N(��P�{������,*�Ŭ<<�*�kJW�E��R�6��x��Ƌ�i��fc��aU�5����� _�]�m7�ӓ�XN��u�e}�������ƚ[~s����6�T���r/e�m#������of�k�	��d0^��g$�wr�n�er���jĉ�`�X�h��[�S�h&����-B@�c�s�I��t}���F���UYl��OZUT����l�ȮX��`�*�սbS��E+pa}���5�Mf�S�Y���;�9J)�ׯ_
��z������*��(�]�4 ;�����L�Ճ�5n�ad��҆����x�n[oڤA�YFrv��������e�~Z�<Y��H�uYRj�(ZJL��(��81�4:c�gj�7!f`s��N?��g�x���sH9N��#�H0�~�{�m�^��c��	J���ox����~�B@{����T�����~��9����/��]l/|>C|F�Xuϒs�z��L���<���ڬ���*k��Z�:�7 �>ٳ�\L�6*Z��pSI-������zђ2S���M�3`J>�.�/��=c_Ζ��G��3d=.�3Y�ሹ��v��Z��4 X�����6�#Pw��0{�A���+��16gƥ~=N�2g��U����JV_r6�(�����,���]��㏙�km�}��C�ƺ~���c�uĨ�Ø̸���uΚ������#���p�	@�ד����KH1�{�ٞ��( a#67g�^g�;+�>�}:#C�4�v�����G�@f댈��!. o䜇CQ���w��P{��	3����������=Sތ�L"��f��&P�e���� �E����&�E�lR\�"��kF֣�h��샒���+��퇅K�<�,���� %�dڑR�쓶޸g���&�6�g�{נu��#�����l�c&�on�9�$�ߒ������u�~`�t�������ju{ξ7��;�g�F��3����j� i����A�f�X��̡�L�b�3�>�0V�C�ْ%ì�������xO^\�v���3ˠ�2!G?({�!$���.-��e��?g$�т����c~{��\Fȉ�=ə��½���Ob�<E�G?��tF��b����2,��Iι���Y@crpb2&ac�Ln�~ �9�r��	���hu��r�s�[,�Ui9�}�~Ԣ���f�ڈ5���ӱ�m���+����g�X�{t��1|G�Y�C~���������1� �!x����_r�9v���e��������&!3�X� �X�+LL��5��}�~�\}o]/˖����j��u��ܴ�]�E��6sl�c�S�ϲ���uԓd��Y����S�E���WR4���T�ջj��z'���3���C�8��sxyy���]H�>{߁����ϗW�����ˏM9{2����	���^0�Jj۾��K@�Kvx��K��f7�9d��� W��Ř"����(��F��cĶ�4���e �Y�قIM����:��%�f���%���j���]W�xHg>�8�������ޑ�B)���޻z�d ��6P'��9 ���\*&�b�뱞��v"ʓ�Nn���{�������lZ���}��D�%�-0蛜�3W�J3(�I� ����FVc�Yj��<+��"�ˑ��۳1�7y�j�������l����V�a.���[w�R������3p�� �|n��u�t��h��q�mb��b[�6j
ĭ�g�'�g8�*oif8=�V�U�ϺvVϪ�i�Y�\+����#��������#�m+v��m�l;�羳y�~�t4���G�h!#�أZY�'D��\)���;#1@�g����\��I���Cq��B���K�~������BL	�}ǾGĸ�eGDI���a�6�y��w@@r���j@ItMJ)��i�FC��GWۗs�}��ܜ�Q�d���ͷ(��B؂g��%P�E�cvT�Q�'�-D��4m����y��E  �m���̖��le��sh>kM,�gc������	���W�xP<VQǌՑ���Y� f�� �f�]�az�:B1CZ�Oe<��ȍ�b}�=^v�������u��W���e]�|ݟ}�������Q{5 Y��3��{�B �v{�ʘճ��]�6���O�4�n�w�9:+��;��}f�cq�Ε��g�w�0b=O�.\�u6gόU*��+�u��͜���g�%I�ٽ���lf�ڋ�(���5�aG��C)��Α�����Hz���5��f��(�e!��љmc�?��2��q��'|'�����#�S�w�j���d,>��9�R�{�������w��i����3���b‴,<����{��j�Ϸ�7��f7���~t}{�Xb�ً���͛�/}�}���<AD���P��ژP��W�[����*j�X7��2����ڐt[�]ܶ��]?ە����u�Zf�ܫ��;�L��o8=�d��+����eu�8*��e����G}������ԇ5='��5cg,╶���O�6���
�깮��l�k�9���[�z��Y��ȱ�m�[Đ�j��;����M�fK����(	!I����ףSC���Ü�_�8�.����s��|�M�8��%����?Z!�����>��\�uRu���8G�g�	+OE�n��Z�@�8o%�%/��~������x��.����N��&���FN�^ya]�M	���� �2�!a�Gkc�mc���pV!]�9��@#��3m?�E����5{���g��B��m�1/g�t�:�}gʘ1VrgvV^��1{��ٳ_�r��[�]o�S��w��n��\�+�{��+pwUd̀�����lv0�ꚍ/	�r�"4��f�����r���sxtޡ�o�[Is��	 e��Κ���_O�5l���}������F���`���1�9{��k�,�)f��JD.y��k:Kv�)̥g����~��r���,$3g���]�^�m/sYဵ��Wɗ�L��~�#���
T��s����<�����dvm����'���%g����������n��s��i-->�73���y)c�Jx4Ԧ	����3�;�LY'�<9p����"�r�������{�97K��r�
�ׅ��X��@��l��7{�nm�o�����/^�6��J393ƺ�0��b��.�,��=3�h�����r�5�V�k�\k3ӀN}��Y{� �p��X S�} �qc��i�~��ϲz~�9f̹Ū[cl�;K��At^���%���gsxV���Ԇ��������Q)&��4��Zx=k�m�q��oAP����O2��Q�kpi���r�+�������!������Ŵ�w�=����Ό��=�H;�D" �o-��]�d*;ڜsmW�T���Yi�Llg΃�ط�/c2;P2r�]g~�4@��(�X(4�L�31��ݢ'��՛}~ܦ�|��70��"�U��l;	4�x��埭~
�C}#O}u��9`���ǀ�=k����g��:7:]�O.���;@������|�A��LG}*ʶ��{J�Nۘ$�`��� ��0��i�����x�����Xmf�HХ�[@�hS����t�4��zk�=����	���s-Ӂ��WV@n�Ό�4�l[f�~����3R��Dћ�8w>�Nڃ[��١F�����7�2�77�p�}R
��k�|.�l>��A\x��aK�w۷�"��<'�e�*^Y���!��&W��H���\eAsBM-	`�Cm�)M�:���7D�_c�)���_I�0�'0��m�15�Õ�X�'猘�J��Mu�דJ��k99e`u��Y{d��uk�����"j�/Z��'@��_3�B����;+ i��*�����|V,���_@/�56ej��j��\��F?�ܰ�� 9�'��j���ׯlF����"�0���}߫	�Y�H�я#o�n]��������ﴕ1��#�b~\�5�,�ן9䴺X�c�Z S�)�>�����ޱm��k�-Q���r�k�q�{��Mvfe�'�-�����R���=*�#R=�SB���ھ���f����.	1�#��D���)�x�k��"�dlS`&��&�d�("RG�>��N��3�ҹ�N��� &�GsN�3�apH�����������E��ǁ̠�@�>c�-���{�b�Ƕy���bA�,Abs0r�s�v�۪��~��2�2 ^O�6SQ�w ��G 8nzg6S�NK�m��e�I�0���"�ml�=�>��iciv�<��o�v���{m��~���������9�u�fƖY���ke��z�g��ʖr&'u_F����fj�Y�$_�c7f1I�j�����W�򳳢��|��;\	�g ���l�<�ѳiteNq���o͑�e*[a˽����0����n��fR���W��U{�wo%���1R#��L;��������o��G�W�J�> ����<������������3"�D98��R(���3�����o	�J<Ș�2����v����6
B�C�n4�m���S �-eW����r*�MX<������{ď?�r�|fVB������^����h����m�W�s@�;r�'f?{����{=��e���zA��1�		 ��z���-lh/Ų�Z1��o�#�iŌ��������ٕ��³,#�F!�~�ih`a�n�>�oV��V��sz>6�� �qL�y(c��wڜ�bW	0E�����������:�/0e�%��ku�Y�$H��F����B׎P� ������,���.�9��E�8�q�@�|�3�9a3ǿN+ �������l0F��!=��C��o����m�Z	}�Z��[�bL�Q<�,.0�SԦY�X:�ݬ�}Zg#��p�����X:ݤ[�����h_@�+�f���=���������;��m�p��KΓH���l8~y!�ڟ���9�zb(���|���/�	���w�����L<����b1+9�lVe2R����{l�x�;ܝ6��n�[��$Ӌ���j�������"��<	�n�*W��P�Q]��P]�[@�gi�����v9�t�{�"�LR���HJIK%sU�zG =+�L���1iG'I��Mڊ��l�6�o�D�a��d�)�N����[ M���5p�`���s'q:<��J�gp���t�4������ˬ�E�)�����>綮����)�������&˰d��.mVw�؜ M6ѕH��ϫ�Qt�2C�>@Y��:wt��n��U��m�׈Y{�r$���	�GW�6�}��L��]�5�Ci�"Ǧ����F8趝�3{�L��n�����,�09xN�E�n΢�Hq��m���ӫ��	�9�<�R������9�L>�I�	���ə^tbv*�!�G� WS���^y���)�qӖ�ϋ�t�v9ɣܨ\|J(-^B◀�����R�O�,���`��3|v�k �\�bgF�3�guF֓-G�1Qs�;�HVBz��4�:2gu���c�f�̈���ϊ�?�wG�)��e��s�0� ������
س0 sVz%@�`q�LR�p�m}�
����� �!�$`<�����G��f��ׇ<>8�iӊ	���+Ƕjph��y�{Z=�6�8�nZ�ՏH7n��z�ys��8����[Ɲw��P��	�S�O~ڰ�{�e{W��s�C���q�c'5����=S��A�F���,l��ma�n��V��1S8%N��z��ɑ�ر��v}ޓ�� }����p�#�Q�����f�$�aٶ�~΀[߻|�8zd>S��_�ڑsB�mєe��k�g�UfXl���"���Y��3�y���v(뾣gz�8�D��mq���Ye�<��cU|���	�oAl�6;�U�GϦ�^�n4��`} �̫n�l�j�Yc�m���֢�m�{���ح�c`r��F��6,�~|�Knmi[�z�����x��k���Y)������'l��`S��*hfX��\�Ȏke3���6뻛|�T��:6��g[�E�!9g S"L����U�#@Y��c�������ߐ��2�rI}Ǜ�<-���gRg��s=U�������3	W6�X����k�n<|�u��dւ�j>x�����ۛ���඼h�pk��Ƅba?�G�
��p�aO{y��t'm$x�Ł���I��Q�t���4~�~v��g{O������V��rٚ)�L�f����׌���Hf�dVY��[y�h�N�A�d���a��]���q�ۧ۬Y�z(�0n��@R�h�][�&����w/˶TΫq��H���<���@��W^+���s��G<�����vI����bπa�J���?X��Rd���i�V���5-�N��ʗ�<K����&��X�~[��c�/�r��t�8n��2ɑ}y����s��>�2��T�w�fR��r!�%��ƫ��|��|����;�$��3$�6�ٶ���sN��cN�b�IQ]8*V��6bI��z�[X�/&� V����!����������:����y{cs�|u���iOǣEI�@;��]�"����I�sBp�'�	e�c�7����h�2${�=;V �#{6&[���@3ۀW����ea��_=��r���������<�g#+L�`�J&�}�����=c'��bЬ�lg�@��١�XP�j�)�w7����+�P;����`�p��X���X�n0�qtuX��gl6���C�����ㄶ�Ǿ��f��$��Nz�˲��zs�~ଁ�8�Ҟ���"��$zB��Z �-�r8w9�/wȑ.���~�|	����0Wc�\�W���K�o�FSL唝��)��|/�F�x����yV,�d2W����j����W���H��i�P9�.��s��|�s�m).K�N�J��kҝ�M�o:����Mh��ݛ�޺G�Aj#�iB̖��8g�Y�-���R�K�,�c�~7�c6vBџ7�@�xg h�>dy�;�S�.���'b�
s9&� �����K��B=��1s��$���;��xv������h��s۴*���@Z��*�X���!�l�9Οv��G��v��,u;��$Zַ���,����� 1�0�ϳ�~=�d@[��{�~��m&������Sq���B@f`Κߴ&�8��wW�LW�1��t!���e;�B�d��������{�D��/:_E���ם����)�l;�pր}����h�i��/� �Xۈ���V��A�h���M��G8�����k��0�a���=�A-���]��FnS�l�|�<ɜp�ޤya�63�,�#�J��H�kl0(yFYW�G��כ�u�k`��_������׿���A昑���X��������k;G������+ӌ�cS�/�y���a*�4��[��W�|���G��9V�93���2s����T�Ϝ�����q� =@¿1��\�wHf�j_����b��Q��O}���lk�?eZ�چRo�r���R�YO\ҟ&_�ޓ�_�7^��(�9��<�G*/��RQ����)�T��[9���@��1�EB�Ae��=�RH��%-�6v������tbP�S�@��+"��(U�܈ra_`,�b{�3Y�"�m)��cs��A����[�� ����_�T�r{�<�z�K��xR@.�����x ȉ�7�6�\N؜�� ݳ4����� �h������?���mۦ���v��6Mt��T6h;�e����e涎���R�l����Z�s^��a��*�$[��@�<�I�eK@j���\����P]'A�����N�u��OR����}�+����e�k-c@�m߶�1g �+ܓ3r*�*���Z0yd�����<�E�Bӱgv&���֜'��sDN%�`��*^�)�A���.9Ҽd���=���ªe|D,hC?~v_�>'�'���e���>3�xvp�4T�'�%�x���=����0��@�yDֶ���4���l�)���W���.�5t_ʹ��%Ţ�oz��u�0c)g���~g��{1S+�3�qBY�G�^^^���/��ǽ�~`�)q.���v���h�S��o'س/�/b27d��v��S���b��)��p�<=�#lb��7��Uh�a�u�����d^8ݮ�ì.}?;�;��6#�X'{��m#�~��.$����K{��q�D3,9g���!lض�1EZ��UQ���;<�8�p]����m{SJ-��E
�I��9 �b�o�� ='#�o׳��3��}�z�tz~;S�;�C�낡=�]����c�ƳT��6|����a��̓��V=�ش�aA��7��� v�9�&��)�B��d{E��B- ��"�׾���| *߯l��`�$�}�~�q��vK�Y�!Z�S�U61����3��nM%&*�5I������-N&��y�n3<���=��J#+���8���� ��l�2���|ߧjrk�1C (/�+KȑQ0��G�I9#�~��D.�F2�j�v2k�`��:�V�O�2���HR9��E�fw�I̛���}���H$[�m�$s��9����5�ɿspnb�����A��:�	�M�T�N����޻�Y�g����gD�0W�#����B�zd3�7����Q����82�z<5��~L�璑�;[���"�\����~��:��F��΋�յ��R꘸��$��9�*�9�1�-�)��4'��띞����|��qd-�;�?��tm]ܯ�'}m=uϭ���U�Xy/���{�9��R*	5���#���3r����x'ӥ�X"-P~u��j���d�*tr(����c~�w�mC/�܆-��B�s7�#�bl�+���P,Og��̹�w ����~ѓu6�ρ��A�S��'�Z����'rdx>�էʴ�3��GD�sfOK�arUZ?6,ېR��8j��R�G��sv�9�0hJ)c�Fo�F�=-��g i�^�X��)�8��:��Jf���?z-���R�&F2�H	�@ӯa��&���8������ ��a~=}O+r�����6�z�z�b{.δ� ����jx�/��c��:��GE��3��HR���X��s�X@P���-�w��=��*%�@'�˃H�zN���ɼ�F02j��׷��1��Q�|���$_2_^��# B\�I�I��O��(����C�<>��m#'��6'ň^mg�G������+��W��r�g�fJ'&�^�z�0�+09R}Xz�VSo޳r�wl��|c�+�v�K�y�7ǉ\���� �@��خ.�l���P���	�����@���3k�I��4ɰ?RE<��:�y�wډE���^�Z%ۨ��mF�#K�Հ���kQK�}1����J���۶aߛ3�уf)��~��z<��}�3�tn3r�=+ y����]���Wt`����|��s2�i�1����,��}׍a�փ�P�
ɘƽce]#:P*���7���-�pُ�&袵�����~���=��% �4-�>u��O�ĸ����3�s�s�8�ijH�SQ>����=�#�d��f�3�9�ʡ��os�R=&p��8�'���a) p(�?����z<;�o-?s����K@�{� {��?_o���HؗG�H�pt�f��o�F�I���,��`��n^��#�-G�*��h���]�T���)SK�\s.,�g����m|���b�>S�GXAi��e5U����)�mA|w�h��$;g�6PKV������$�Ѕ�9[����Z��r�H`T���l���ʧ�-�[�m�þp���]���1y�'g�9+3;��]�ٮ��LE���ڿ����f��3σ��(!BJ�D�Z�s��<:���c0mȻ��g�$d�zMۉ��2���z���ֶ�J��R3�)#^fI���ӎ8�k �j�4���C��:�X���5���9���+c����rm�ܵ�
����K@�?�{ R�L{����=�j��2(t��g�[yZ��3�k'��sx�=jat.��_)�����]���}�~�a?�dY�<�G�s�A�6T���\5�?	�Y�g�&�����:f��eȟV9��G�40�Q@Ăo2�)�9��@%�׬����	�M�ߐ��.��!��I��
�zowf�9ufS��������}a�����G�c+︼NV�_h�m�T��� ��G�a�j�є'�կGq#����&ƥ%m]�qWʿ`��R��3G>�5�4��w��S?Sf+��VaA�ip�����r��Ԥ���#��s�iN`�ŗ�lB�w~oR�]�k���/w��;^���7x$����`�Iv��Ϩ�SN�Ր�Q�ח��{I�r}2^���;5�OT�[8��;ɬ6��l��Ex]�Őro�R��5+O}ޑѽd�9^�b,��G���Eߊi�m�Ɗ7V����u����6��|��K`�ʼn~�z�[��^�{�c��*�W�L���8�ǫ\�3��n��M@-��y}�!��߈����%0b�z�9��u�� ό~�}�#��lq�dHz�k�?��^n�\�����< Zc�c�=�*��g�쒢�Jr��YL	�%=1���`������� UEXv����@��m1 � J�^�"5r΃C�l~�8�j$j���K�wk?�����'_^^h��;v����֮gM���3�K_���k
�Ŭe.�G��K@���������l��� d��Q��m�d̎��	6Sh�`,�Z�&��~���;�������j�b�� ��v?���%Yml�E=Y
frX(T����~q�@��V�w��.���OL�D�D��eR�ݗM����y����;������­2�I�Ѫ���XG�T@����c|T�9G��|X@Gہ�T�2����s��U�i�#�Q��%������YV�m����ʒ ֍���6��˔�R�:�ڡ�b�lk&�9�?~�5�b�r�t_h��<@o`ڹ�l^�8��}+��Wm�A�[�d1���z{{+�*U����32q���9�0ReG��t�'OZ�"Ꮯ ƈ}�k�Wm�A�ۏ���������{/l#Kx.#�Zo�]�H��bs<`���RwL��Gm������d�CSz>��0��� dW�O��}�8���Us�?I"����ޚye[$�#�s���@�yMu�J���~�w�z�sa�xۻ�3h?��N���Ә�4fY��tfG{��f4��om��ʞ�V$u|��3}d�Et����ϕ/���������p����e������t��4�1��������w���	��6b��E�fm���A/�`W5�\܍�Z�V~DX��m�=�UfP��7�cq����O���梅�h�~ڡi%=�A��?;b�t����|.mΩ��f�g�����֠~^���6��9�[�#�h;M���d7��9~j���G���Zn��d��u�@����?�'�,A���:��z ���Z� ��r���3�0K ���ۭ2�Vټ`��|$@{ ����R��,T�˛�t���Ɩ�����_t�^{�<`н����0Ve��I�I�4]�T��5���S�/�S2j��6�\/�\��ϖ:�S�{|����hι�O��Q>,��_ng��e8���
��5�ˌ�R�#Cǲ�n�% ���������;�9!��g��:����U�'[�=1�6|�9Llpt�zk��iZ�d���<K+�1�PKȖ�	2�j��^���>8��(�ⶡ���z�yY���`N	p�mLH�ǫ���N���b�������d�Z6����[�vpZ���3������&G@��<���ͮ�� g:t�YI�D��;f{����~4�t
�GD�b\Ҵ�Yo�N���:_�A��>&u`�rK����|	ɚ�!C�kD81��\sz��N�-����t�Ve�L�I4��&5�%M�Dk�6e��C��#���k{�5k����J�;�?}��8��x�#����?������g��U6����6�:&����F9�-u�J�;�7��+�A��d@�䤊8�:��MO\H$�x־HښƜ����*{��1�\%eMR^�y�� ����i�F������*��N��:�2�M=o���U���\H�ݽݝ+����RW��ަ��W����ԝ�F��nl��a���ׯr=�K��-����~�7�����Ǒ|O��#7^m��k6�ڱ�s_�,;U���o&����o�b�*{�^Gc�lsn�Ĕ������Уd�)EKu�hk�Պ)���kU��lc��V¡�|��սS����!WE?�s�ƠMU����w�����L��ǈ�W/�>�����|	Ȍ{�C@���K+�@y��n�)����P+�y_2t��4R��2a\�T(��i�L�h��Q�c%]��"� -�E���[��Su��gnh_3�?��I@�@E��to7�^��m*�ɟN��j���9��e]��仌$*p:�4�O��������2^k�<�������+6�}	�M.T ��I��f�{�D��b���aCJc���f����eR)��`������p�2���w�Fn�///�}2�<`3Z>%��9�ׯ_�9#��z���6�u�}/ǣe|F��Z�r�Ⱦm�Z+��� ;R��:�'����Ic���iq2�n�d�s��=�k�X͙�[�@��Su��{�P �nq�ڔr�&��,Y[te����f�mM��x�����i��⛮��w��db-� 4��z�r]�Y���T{�rM�9\b4�`K���Ϥ�ޙ��v���2F*��v#��%��`663�u;sڟ���5L�����+�����|��K�u�z�'LVjt��4RHp)":�zY�0`�g/!'`�T��O2Mr��S?����}�D1����MH�٤1ҀG1��D���B)�ε�b���`��K��q�8k��E�7Im�"/qzG�����gk�0{j�����{ګi#��������	d���f`_��SI!P�u;��rd��s9Գ���gVg��CS?��4峄m}-� �E����}�]u|Qyɵ��1AsS�`6�)�楩��2+pg0�qdG0��~���<��C@Q��h�%�.0��á�73��N2���VRn�����p��z ߱�����H�9�	2 �>��o�b�3~�p	�Mќi�'7X�\UK\�Sɧ����SG ��L�GD̙:\��3b�HP�7e5��F�y,>� y�y�~X��7[��H�ޏHT^�}:�/��}�j���\����4<'����y%����74Op���}4:�P{�w�ޜ��x�V��w���j����ܴ�?F(�6��]l������W�7 "�<��+���E�߳�<o���yI�<s��CۀJ�'�Nw?�{Dڴ9�D�a��ϫ~?z/t0��v�6�� ���1[��6��cO�R�kΓ��\� 3�h���^�я��k{N��°����^a��3�!�ȡ��\/�_��L�8���B���������,�C�)Åˤ
��k6�x
 �o���d6��l,)wz�����,]��#�iب �+ꀕ0��KG��ܲ#Y���g�@�6��W�C��Y�2�����Oծ��q���]QH�;������Ը� }&Y���gG	n�L,�r�>�=#���������5�t�3֕��u�ٶm�a+�x�ٖ����$?�:������1G��`s�j��}߻�<�Oף�MK��J[Cy7����h����Q��k��u*Ձ�s����r6�ic5D�Lϋ����V*���5����5d��8�:V�Gʤٓ{PGP���-z_��st��}��/�6K��h�@�Һ��p����g�����~OeN�d"ռ�\nkټ;�� ����.lؽ����&��@9b��%�P���B���B'.�m���B�b�ivD�K���3���m�|J��/�ҡ�����#�i�y+�ȕ5�[<�v�jቘe�/z5�⃊�b����\O�LU�2R��\�%�����P��zFr���1) �ﱜ�X�͋� GJ�p��2R��K�����V�l���b�_"m�����=�ޫr�s�<&���4nx�uI���#�w@��~��ΖBr	ԍ�4�>{ "7�� �!"��2F@����c�y�쨼�����n��$�"�&��/�wX8ޣ�y��4�-�d5�<�e�REl�b��{`���I�)�O�D_�+��S�;���[��C,#�t�Q�%���C�{-��5��˫�nTZY��o���1��l �SL5�ۊɣ��2XK��f��$�E�6@i����t&�k*ent��\ګ5 1wjnm�h��#S�u���N����9����s2=��,])E����t�>���A�	e]p�6V��J����8W�>8�G��d�����:��Lv�h�ŁO2�F}N,���ʗ�L ]JI�+E����ŔI��'���)|�@q��x��E��tr�ɚ��g�K/��EI��~�t��3��|�"O��)zt9z�=�DZ$�\��نƘ��*�' �:�%�)�Ů��-�Ǡz�t p��8f���Xm����W5��je�C+��41R�]�c���4l�L��3�!��+�ݔ�w4�Y������q�Q����Z�@3к���������,"@��d6�Y����֑r��]X'W�=������l��TyԆɳ����OPW$�$H��c�.��_����ߐ�^!?ri'e�c,7��/���K�dR��.SD�3F��U��#q�v��~���8u�G�ݵ�UB�ڢ��| ��ɉ��8s�T��52��Q�z[�D-R�������5�B�{,;�|*���e��wdX�j6�v����*��]�J�v$��'~'�gwQ�3��Xx���>t _�'}O{�k9�ޅs�d�Ħ����B@�+s64��m[��\�L;�Z}�nϠCi=�p>�����
�Ĝ���$?@.ZU�T�^Jnq-��ꑘ�33���;f�d`��C�R)Z�v$H8����� ?	`�~�rD ~2�8���k��ηLvM��뼔�ˎ�6� �5��W���?v6�9���T�R~�Kp��B��?��|.{Ѳ	Fu�M���|;�:�9�c�"��%;��p����s��bܩ��(��� �="��R��}]9Rm��B醿�$(}2����|"o"��Jv|�(�ˍ%�%�G[�d�vR�ezBޯ�������Jf	"t�m�� ��g�`[x%Y��~��v����������
;2�506��"��C�����/LOq$��Ҵ�W��׳moo�ɾx(�MN���ng�ĺIP�RP���� <ux)j��c��������O�+������7��ǯ^����@Y�f^͕#�󪌱�e%�!��޾����&�1�^�y�����X�� �ʒ`U������c�E���}%��}	UߗA�Ա'�� ��0�ݛ�}�ߵ���u[���^ݧ�r� ���'��7����o�� t�qj��=�.�5�寯��na;q̖�{�/Ҽ�;��"�:5_�T��oW�Q�Lb0��������@���URU�\��D�I��I����gh[n��p-ћ�w��+���➰��5.(�N��%{���9P��H �����;�gɶ�cΙr��wϛYm�'E��Sz�]Le���}�9�� ma��� ��T���m���Jf��j�;�]=����]����BRk"d�= S��#��,��b0���i![�?��E�Z��=���j�ߵ<v$�Nb�؞׳��R�� u��i�?��U̷6>���3��?Y��)D?��O���22�1�1�{�}�~���:�r]��T�<?�6QX�TYq�>��;���K�'@X{F��$��U���e��|x���s���c��T�؞3Rj��]�����~��M�~��^"�}�����F�bD��2����P�?[�d�w��O����@H����G��'�S�+��k�`��M~$ �E׃�P���j��
@r]һϪ�@��Z@�ڰ�\�1����H���H�K	z��������bę��TS��y��C��ٟ9��6�I�<�y,.f_����P��� �B��4�
�sF�DU���-�`����Ѽc��C���]#�1��Y������a�z4�(��=���8:��� �c;ƾ� ]�d{$���a��ڬ�Z-�6G��/mP}A&2�4��u:uiU�ϫ��j{�e��3�������2}X6H�������.I��0��T��ob+�!KUic�g��8��g���~���L1���l6�1�%�?ƈbtٙ����Ɉ _%_��'%ĴW�i:t�G����)[�#p�7�n#�U�ы�v���`���d4ũ�U�5��.d��g��3����pC]�~k��m�=Cq|���N�<��J�Ue�3Ĵ��%CS�s<L�@F���\��v���O�G@W�$�6����==������:�$��ԍ��'�$�^ͼZ��3�4����K��FX(~o�u�T���e��h��Ƣ+�p��Շ2���b�\KGH$A�h���~�%k3w�?�9�Kx.7q\Z=��|�i���.����d��<3�z�G�3�:~�+`���׽���j���Oi�D�B2�E�)���=�u���qggEƸ�r.���a�gȗ��S	*m���tQ8�)��a�*@���߼ʍZ�cJ���\8�@�E����V�װj�d����g-��J�E/(���WĜ��w�5�����N���;c��i����#�sүٝD65�eOj	�G`k�12��&��?��B"��#�}U��y"�N��U���a�i��?@π���c��G7�����0I��7����7P �	S���:f(�������gq�*���'[f��~oέ�_���b��6��[�t��Z�#<��",\g_���kϖ��fm�.}8�}g�M��t�}����Cmg,sǷ0PJ�ަ
4�s\i�w�7����T�U��\����'rfc���'��0E���qtL���;��S����6Ɣ>�Z�.��3���9�s��2O�����K@����~��=��@�ޕ���-'�hv�bQ�*��W*�OzI��K��\J|N�0Hq�YW�&���H�|��J�CvTƳHe%dVa͆��:P|Q�D�qB�\�4%��x��q�ݵ2���V����W��{= ����'�n�u��9�Ǐ���W��� ���r^����+fq�Ƴm�9ǭh}:��bT���^G{N>,�:�9cV����@�X]����Lm��ױ|��ܦV�v�۸�gx��`WGm+��샇�+�L���Ȝ/�4$}ח�hY�9����Y�z )C��Z׳��� �{�KV�{�m{��G�Ì�@�n�!�8�p>���wl\ >8l�[)/"�6G�^�{����|TVA��^��pyOy"Sk
���I� ~,��0y�Z�4� �:��y^׶y�M6�15��ZbL]0�̓G�e��,l�k�5L�|���F��� p��z�0���mn��9��n��t�;�a x�Pv�%d� ���7��f�D��>����U�S�W����<�������������Y�/��ӹ����:�P�>V��I�cgpM�p4Qu]�mZ�����k�`d�ݶЫ��>$P����lP@[l���^t�(�m2�F �hELQ@�>�|�b$�󎜵  �j* ʑAWN�3�U�%���n���жwټp�=ڮqU�sma�fc���~�6���l��<v��Eў~C��mH���q�
�	��V���K�R�!3%�,���l[]��2�f� )�9;tc{�^܃x?�r!����i���d�c]��fp�u�������xh�m��2��~}&�S�D1��l����:_i����Ws�G��;v`N�o��6��1��beY�|���Q����^+��̣�v"q\�n>���gG�To�t����r9Hr:����4����B٠�O��!u��7���6O<	2��8�}��J�3O>�@�Z���;a.Ӱ]X �ÒŌJ�<���6 ���P_��
��NcY���T���~>��m�x�
R�&�]Z��ڌg���~�\�����nfO�RjJ7��c�{�Ì!��
�e�jm>�B����q*�L5j�H�9h璫�Y�ZFf#g��V��YMf0����Su:��_���Srk[^�M$��A���վ/�s{�YYy�[{�.��-v��ǇQG�<���Y[]��=Ŏ��?g94!~>J2�!��xT׭�Ӫ�>��1��O�Z�ږ����{�����	�H%�C�mxͯ���?��$SD���craH9c[�5�|	Ȥ�o�8}'��>It�ĳb�Eh�'Ve��R�,'-^M�v� �s0U�r�)�i��Gee�i���`�{	���Æۍ�^�-���E ��������Ph³Hu�s8L�&�k�:H����A��[��1D4u|Xj��x^hg�+���EX��;�n���3�ڈ��?#;���;�Q��k�,�^�޷�����:-G3�	!��i�Ё�9�W���m���{�ԝ�\�ky��6�n �]z� ��h;n�lX��w6��U�Q}oՑ�������;}���� �*�����M3q���.��7���g�\�. U�1	0��������Y۴H��~���ɑ�~��z�2υ$��$�%_2�� ��n7
�Y,�3ΰ�),���1��&��욊����Z�I�9�1��F4�_�������-l*�%��g�B�ݛ��P����LFV�>�#�e-� �-��Ӡύ��Zn%m�QR�}�X����1%��7䜱�n-����LةU5e�Km*f<����|��yH>�*h�~N-�Y�\90W�J�V�Z�Y�Vf�X�G�i|f�;<�*+)ڥYei����r>%h%���^�����q8Ӏ�շ�m�]	�~����s��86(�59Ԥr�x��Q#}5�]�ȏ6mk�ːJM��w�2������A�|�����\@;����S>�̪%�t��mP�*���۪M�f���.�
+t!�IW��r�him;��@t�~�p���� `����{�.��)ƶ\7�x�@z&52K`��b�=(5��h�%_'�V�\.���+��f˾��6Tyʝ:`�<��l�R���,�i����L>��ރŹ�z�L:�K'I�\�n�	�o��b	�+�Y	�ک0-U�RV`tv����uX�)�ڰm�NȚy��&2z}��y���x�O������(���a�MJn�g�ٳML&���V�k�w� �a _K�j�QjZ;G�K��`����=~>>0�?�u�6�6k�����2�Տ�Ly�AP~�����`���6��r��ɩy���i��3q���Kr�3d���{�6���;�g`�,�%l���Gx�ĉ}��'�B�V�,�r����G�d2�M��g>Cph��#&�\�T,,�$|�Ҵ��fp_mXT@��d�DP/�:qSR��� ]�}]
��^�`������o����b�ˉ�b=g��jJ̔�p0���lWrt��|h�@*�Qؚ�W�w��+1������l[v�=�r=o��Hֆ���{�k�E�\7�Ĝ���Av|t�f�u[��� Foŀ�Uӫ�-�f;y���*3L��#�`x��Ԯn�Dӽg ��S``x�_u<���K��'E�ә��������-�T�r�?4w�9�I������,L��Eև��H:K������!�*3�B�C�|b��}m���1��]%2���� P��x�������<%N�}(��"JF��7���|���d2�$&J�&a�Y�����������U�
����2�'�Ge��foo��ζ�w�\`bܛs��"p.���y7�_o��A XoN�� ���Y]��k����ROɝ�7&+�g��:��0���ݏ��X��|Ke}��OǓ͹���`�B�����xv���8~�l*���~�L�=Շp�R�{V䵫�����ڳ�9�1�g� �&
y�P��|�9aߥ3@�Qf��u�n��Y^L���:����yE�Cԛ��jp#�f3��O�c"��'y��S��g�xk,����{�ZWj]�kUD�9���Q%��53�6���3ү;�g �jr<���MX�A���|�AY'B7x9
~�C65[Lf�N�����9�=7s��r]��������o~�e���i���c���S��~w��01����s��#�+vY=��G3�2&g{�>O,߅���,�f�^�k��R��b��l�g`�jv�X�6��q�vCz7U��&��EV{�Ϭ�;��u��O�Q�(6�\�L�1�$G��k�֟�<䗇��I;���� #��?��j�\g��3�+��6��k����2|�כ���l�]���d�#�fQnQ�T0�Y������ҏ�b���H坃c�_� "���_����Q��T�!Úz*��j�)
$v�V��ʖk��~�լz�x�lw��CTׇ��b����#�R�9XΙԩ�����5k Y�Wh-ٌ�L��i�Q;+���`w6�_�Gr�	O �_����P�v5�k�#��xSٟ�`��ɾ9{��x3�lKqr���	���9��a���AZ����C-ި�C��M��&��5+p�E��/*�,
�z\�4(�uZK	�2�������K}6;��f6�t��)�!�f�M9Ѣ���<��H[;9>tlҸ�����%��?��d�U��Y�ӫ2� ��2| 7����~e�j�k�;7/ 0#��~��*���^��e[�د�Dh�8໱����o��u���lH+}����Yt�3&�鸠��9DU�>��~���c�\mAg�JփWsKյQOW�Az�v��y�9�tL�1Td��������ޜ3e,wW.@�3i(�]�߉⥦�B�u�aX3G�e_�zXG����˸�)�d�n�)D��'���Oi�J��ɤl���Ԥ���F�\������E�|�~��W/�#bH� �t>Z�,ц����&��F�WE^U׬<Z� P�?^_?�Iu2�F�GL�1t��I�v�BlL�%�^�i͈um.�^�i�q;��X�6��B (�r���x���K��ں�+��Zv6�lO���D�iH�♼�9�2;�l<�����pW�5r���ʺ��n�-�[��x>�^�)y�l��,'K�����K3�Ҧ�˶�� �P�Ru�?T!�>j������b�Q�!&��g�+�\UAK�{��y���2��X�S�s��>�w�ف⼃B���s�d�9���!5�w�/b2�aO� O9��m���SHK˗�:����*�aL$�ms&[����'�2H5:��F :zn�v0��<qY�\˃Q�(���4�j��G�nɐ]��v��v#�v��6����YY�֣6��L���@����LG2�dme6���j��ݻ�^�&��T���6l\g�2ϘyJkMG�c��A\��ri;��{ݔ��?����.C�9�)E�1��E���Z۞��>��2�����=��5���<7�Ϯ!2!G���p�sB�n����Җ+eHbE/�iO+8�}
Z��cT�v&1��%e/������r,�;�~G��'��=�h�d��Ε���_[����f�>�:��w�v}�e%��/���頖���(��J�߁>�k�����I�����F�\�J��^#��?���������N?�g�>��7��T�}�����+��(�S=5�,�Nn�-��<�'�ȧ-3\�u��� �.�EK�km �2�#���}+CY�M)S)&�{Ķ1Ns��=V�u�J5Р�/eD��$p�Z�^Xc�Tg6'	�,u��{s��}�������@ke[�����yw�p�����H��,&7ΠRBʘ����b��m�w�����i!��$����x�R�^�t�B�̹��U?�g�� �`N�ӾҎ�Ǚ�K�Z�sY?���(��I��X� �g��Ld&���r�fB`�|܏<�������8[O������~��9U�C/���[m�#R��9�F��8��rInq���˿mېr�c��2ۆ�m@̙�6�}�R���h���i�b�w)&��3y�֓V�>g*�=�L����+�d��c�B���g��s�ڈ~�ߗ���o�N�;��(�x�޷lFGv6C�B���BɈ&u�����!??R�3 �ކGl��<#�{:��I1�l�ZkQ�&R�ӫaUV���$վ2�9@�hya>��j�.;�N?�[ZϦ�^�o����=p���Zx��	]3!2��#��eR x�^�� bW��Gj������|V; tD�p]��#VO�[�} #W�
��=���A8���:LW�oK�����]�H�L���-��f(Qe|>w��(#�H�_¬�YM�l)��,��m2�/� ���Rxl���Ƀ"��*edO'7��;����W���Oaz��"M(���a�훼1�֋Tg�1U�3����>���2���|�I���>��J��e����[�e~�XL8���jG��������M\���a��Z�ʶ��n~�L>��:��2%pw�ic8|Zض�eV��=�Ye���~�Y.�~Jo��s,}�|t��fV@[�Yr�,��ð��'�+��1����ow��紜u��˹�XWv� bwȍF|��d�]M��n߹u��k@���*�孎��!?���~�|&�"�f�\=1w�<�Ģ,U�G�9��m�%������ڵE�d��VgS9���7��y!o�H�ν��H��Km����b��TL$�(�u9|�^� I�+�,�%����1�X~^��Bm�Gu��	�YEŲ�$��Yɕ:֞3by+[��6i��3��	���~�k�Kk��Z�]3�)�°�ΞP��>������]5Y�F�p{L�{�jV�1%�mӄg��<g3�Ȱ�T�u\�U�T�P�?�3�?��;I^x6+d�mHk��]?�r�g|�����Ќ=y�ٙi$���J��'�b�aWb��1�%�;�s�@`�@Y��$��+��ns����~��/��y��o����1v)����y$d��X#9:$W�<VpI ﾿��� �	Bo �����܊q�w�֨�,��仉�����g�z___���l�r�l5S��۵#����Ԏ���k{֔@�Hv��`o�����)�[�r�$l3�Q�u2��YՇ�lI��g�Jz;�ƣ%�w,3��M��c�L�;�#[���	����U*k\���d����Ɇh�5�l�� umm��ޜ�z���i_�	��r��S)�!B�d�flվ�e:�}�����Z�o�� \yFG�!���|d���h���\��=sb�4������X�>&�0��2&%K�>-���x�����"�{#d}��!?��@������ח1Α�sG|��Hu�4H�8���Y�5%�|���{��|͉�����-�+f r�J6�#V��d`@BJ�{�yM��#9҂�����7���t�#Œe���QR��5%�&�3�xyy��~/��)�O�!lۆ��c��)���ƃ�w�/�aaC���W��Na %�%�I�V���a�A��.%���n�`$��G�{��'��o_����k��<k=���ڬ�C��]q[���Ru����n���oM�W�5��
��w�k5� g77Ї��H���7s�!��1����V?}iͦ�U��#�_��PhfR&�W���4��,D%>{���_�+�(�v�!��V�S�/Ie`����5He'M::u�2�\;��q<TBdЉ��Jzח��p�u�a���ck7��)hL4�O�e����d+���V����Z��)浟2���:�I�u	l���	�q�[��-�v*6�ۊ�D��۬���˲�u$W�Bo�v�u���ߠDf�H-M�ͷ7.�B�j���#yɘ��SSK�@�_"���'g����kw�/�Y�`��1(��)~y"����zG���m0����m�����ɂ�-.r���bņX��������b��c3K�c��-Ċ|B׫���p]���*Z���X�Of���&��Ql�,O�x�k�w�(v����z#�Q�=U�~����>�O�pĦ�{틵�I�E��;бH&�[q��Q74۹>P����4�-���X
��p3�}�� ߐ�ۯ7�|^-�g��f{��!P��ښj.6{ط�/�n��4Y0��u�:���Ҡ��+$�tܼP�����з,r%��Q�}3���T�GϠ�ۣ�f�^�`;�/Xu@�d�ɇ��gH���^��[�u��-��	��5��ϥ��5���K$�Y"��k�M&�>�d���hWV��}��:�jgR�+q�������;PSa`s�.&T��LfV��1"O�<ó@���ܤw�b�i_����DA֚��h�Ys����"v�3���%�%Va&��pAnT�}�g��-�_�~�`!�s���q.g�k!�M��IH�}�;.��.I�v���?_�T��-�~w���[�r��Ȧ]$x�VI���%�����x%8K��65�6q�����D��jr١8�,K��w��;t��Yn{Mgh��y�cuv�
�?:�K�����O��Ä��17T����r�v]��`3�R(�?�����8��!7�7���vH��j��t�9�9��z֌X��x0.�_4(&�s��e_��L����Hk����5��oɕ����R󿁊Њ�{�8n�'���8+�6�!Yǉ)��H�0�mFbڮ��w }�L��v8l�`��8�̝1�2� ���͍ 8���z�}^�Q�aU����g��Ͳ��=~Qg_���?��!��z�B�즠��X��S��M��Cl'����kX���}Q�4*a=q�~�1�ӭ:0}�C�|�[�M[�{~�|�E��XZ�� ��W��՛���ed;?M�o�~ip}8��L>�g�$��B���D��������I�ˌ�kD7����~W4�G:�%����S"��G�)T����Y>�s|@2ŏ�M�ϳ˨ب��'7C{��pj�Dt��k��6��͊�Z��l����ț��B�j;>K�~yB�
=�t��U�nmOP��-����a�r2��Ǡ[��8�c��֪njؔy4"�5����~2�M�R���Ǫ&�K�ƀ�&�a9���ÌQ�r�^����'Rj���
�jˏ`���d�8N�>g�W7�wT��{s�n�l�m���#�3	�����'*q[V�NK2�������$m����59"���.��rrbU��_�(��ZNp�l�u������m�=,e�/ֲ.(*r��[t�:��JB�)�8ADA1��T]�~dNoX��d�~;�M4T=`2� t�_M�0�n=T�c[���6�Ӈ(�Iv�����m�	\�>5]�{�#<�˯�s2���>��_�h�w����*�~�+W���F���b�3��u���d~����ښg��(��f���P�/tB�<,՗|�5g�>
ݺ�C����.?�_j�.����M~k�h������E�S�;���PU��f9�Տ�O_(ڌ�K�s�������d�- �%�Ys��X��xqE��ve�D��0�!��3L͚F��p�9�h��Com��.J�\>��X���g�_	���vWc�љ�=p� 7��C<W��~#���v�6���^t���%BJ&�ߣ���ϫ�~I2R����հ6�lY0ߏ�A}�rPk���_E*18�>Eq�<[�K����:+�?	��>WD�wQ����VF���RpIbcl�'#��I�z�%?�r�迎V�S�w�5�}ъ�-~q[~�9�����W�����y����0\Se��wd��W$<��o_�<Ώ�|��V������Ū�;�4��������$HRy��φ���\-�n|�"�d�(
�ҧԨ��2p°	�=���l�f�pU̾:U^!��Y���vP�D*,F�é��eF�FJ�r'�Ŧ�;��ܔK����M�ȱk�����B�0��<|#��|Mf�k�e��	W��0�uۡ�}���XTL)��6$�T���7B�%$�Nc
K��x�C�/ܶ�;��'�+bh�-Fg��ӝ�߆���0��G�{2lY��E�Ѵχ�Vd��#���[����[��i�@��c��i��fן�[ɫ�/fO�f�AJ�j!g�g7�?3U��!3�X^�x�Ihmlߠ��W_��D�ֽ�F�V��?���ǝu��ru>���qJ�v{�@js���jVj���Z��cj�n+����e#t���LND`39L��%g�F�{�mC�p�z����a�\v
�k_62�ȵ�FxkCW���덢91Z[+
��?"
>��2��]�W���g�)�SWWx����p���NhTZ�Rgz�'��o�_���&&2�e(<�&��S�Ӧ����$8ܲ�9jTo4ש8J]�å��҉��k���NU�U��@?�ʆ�����5���U��r���%��F����)P�9�E陽,�0��n�j���
�֗HJ�}He��9�+?��� h� ���� G$c�싅I�߶��6�g7+����E��ѫ�voF�٭�c������?��$��z��P���gK5j��1���3��:Un���n�x'W�� ����(��I�� +��z7�'?8JWm��5*8�T�_=Ų����� �R���qْ�T�����ۣ�&r�"Fc�
?p���5��{u�F���M�X��$|cY,/��NCAf���L�aU83ɺ|�L��1!U=�z�[��>j#���ȧ�u�N����ӷ�^GU�"� ؙ%ƹ�~C	"����S-��P����d�o��M��7�a�
W�n��&�z�eC�R������_2J�g�R��O�c�C�G���gbb�=�j�H�����,q�$�P�?���e�gL�J@��l垎���Y� �M�w���Z�51/����6��Y�J��T����
㸄�3�9���� �������)��;-���J���g�<����.�0ES\q�c>۶�ΞO��p$n����H1��q}W(�~g"�=h����S�Ӵ�ؔ�*%hm��#�H�-kz./�$�)�3����S%�.)y�uy愍���"[O5|�[P������0"m��S�y6��Ⱦ�B��{�Y9�Xu�ζr�`QF�z�ݶ���<�S8xʹ	��&:���x����?����f#wv��!f/G��;�[��4��5:�(�zIp�O 5G܂Ӯ%o���e9�$��ιܣ\ZL�}�, �
9��� ~�̙où,Г3�q� ����X&��vj�h�x�v�g2E�q�u��6���U@�G u���7U� }�	*zސ.A�о��X�@�,iM�<i�ηL^&��h,���_�Gs�3�D�%�[�/%��c[ʑN���v��&{�h ��:���
�S[@;!˽eOs馍�՚�W:���k�	�d�:����r�n�;���j	~��7O�z$����r�Ry�H�j�T��l�~�� \\F��`�!�o�9�^�\�oD�F���1	�$һw?h��l7����dZKj:�L;5�'7�ZQ���7p�-9U�l�A�RH��yf6`^�Y����<H��z�����e�p��6�8L7L���L��*���.ӆٻK�n��/�oy��[�$��wo�hfGlk��*I)��-e����d�����2�1+j-gd� �	��Fܼ����kZ�1X����tZ>������"y6����ݷ]}���ep4�[]q�!_c�?f��G�;�hZ6"~�/g��϶��m,��u=��U�- x�i�g�����Mo� !!�|���}X �em��"O�3iW��9M�8���d_�n�y�D�dt��à�ikg�<P6=-g`��"�O��?�_]ybA(f묥�$>�#�B9��׮����0)��?��1�!B�˟g\�;������WJ�mJn���<!s�BD��X��f���*g��PgԌ��Ճ�e�R-+���°5mDP�[PY.g���(Aݿ�������=�	��}�Q���5?n�ܠ�U�2tC+�D�2J�dH�Dƪ��;����=,p��{��͈ᝤ��7�B��c�׎-a�W�&Sڰϊ<Dk�aߡӞ�����9)��܉n���τN�|b��%<&֥U.��F�_�~)�]dÆz�P��q�V�9�*�x�����/r�X���4�g�����3�_q����)%.i�-5��)����X5���j���� ͏v�K����Txb���8��h��\��3���f+(O@+��_[����*@Wc\�;�Mxq׺o�l>֟���7ȶ\,��|I���E�d�:���ui���;��? �&��K��'�`�r��&ۢ�n'u)^I���&X�?0DF��d(�����4��^�jk�4d��П�b�9�3c��Y�:�U���c�!�఻9�$�Vsw��������"����F~r���-�7��;�[��&�b�>usOc�M�yk�����[�d��G����[s���h�.��6  �o�i���)ys�1y�Hn����]����\��޻�O�b��

*MП��G���L:�ߤ�Ok\RF�Z�~��� u�ZѢX<*#ێzєZI�<�j���؏>�0[7l�Q[�i`{!���wu�nyO�X��g���c���W둗�"IB�������p�vKE�e70���i�����x�����֋V�S��ui�3�5��`�T2�M�ۤ��?�)m@�Ŧ��߿W6���v��� ޷��}7��*����qÃ���3K۳VT}3�'n��&����"�Cм��c��6¯Pф��'���#��L�˲Go:�D���?��aku��*ܿ $��y���`,Vh��f��E������욞U�{sYO��w>���� z�͔a��~�j��<_dS�H�Jo�Ĉ���*.�#M i��l_��n����}׮n;��DN��ff�� Q���@�H�i�:�W<�g��B:
����>��F=k��˴��!�<y�5}
G����2�`&u��������\M�Sq��N.��I�35�sG1���`�p�A�A�չ�����]}M�ܫ����{\ͺ"�<����/�w1޷揗a��>cu��j�����:L���K��k�X��d�a8RL�g	���B�4���v>:�ݖ*d�>dm�_	QYC�r����w���=��cT�[� s��;�P��Й�m��.'��y!Ca�h�;�]�(���7B��<�@�:2����i���xy��<�e2^l/�Ӱn��Ӹ:��Tw�j��P���u˺U�:w�J��ώ����Jg�`vyv�����v�fH) =�k���Ogѯ�}�`d�{Ƃ��cb:�X����yX	F�3|����/:�L7+��Y`�j��{:�:'zq�.r �1��	�P��3Q��)�]޼Cq-�u�8��;Ki�e@{��TK�X-Ʋ�M��X��m[����UC�#���Z!��(G�m>f{�4���>�<[����*�Ǜv�Ӂ��w�������kS^t��	�,�;���]�xK*5��;G�7�l������9�����\&�'�ĸ-����D�)�z�f~W��U8��v�i�2�x�Pq���]�y������Չ���C��ß_�5���['"j�Vo���O=���� �^)׷Z�F�%^�$:�)#>�֚����59|��6+q�� (Ղ�4d8��"٘�UH��y�	.�KA�y���Y�e3�D��1�0�\.U���L���x�Rԕ���rEI5��H�S�V��r���B��s\�je��� �F?�x�&U'�� {EY�lĩvk��i�ߕ�=�z�QRU�Gb�aΉ�d��f��#xqlI��ĵ�!��1���[��ٙ��/��D�k������2��r�,�~Ws(�ٓ��i�M���콹����P_� )s��Ę娜�7���qߜ`���LEf^���s�/��^�*|�]���**�R��qq���ef��p���k3�b��$S��K��E>Z�6��7FZЭ��7�����U�T���P���fW��NHJ��0G1��>��]íB��C^�P�^nW�U��*�ljf����#�&��y��䇱^?e�7͛�>�x��l�Qە�S #'_�̅�jĜ�[QգW�Q�l���9��mÒ/�>����:�y�1sVP��3&A#����Y�L� �V�c��-��v�]6]������'�,;����49����-9J��Rz�wj5��_ޕ�K��m�󻞮�(��n�d�xK�}�rA�~�T�hNd��M�+�i[N�������B>�qQ�8ѫ8�k��ӐgG&T��\����%G(���dX�A�45:�^c�{���)8.���'JnPW
���w�|��O��e��/Z]k��^I��YD��2�FN?��N�U��=�ҍ!��ጙ���Q=��(<>w҄���\�����C��Ӱ_�-����[�iY,���b|��t\W�N2t��tZˉ�2U�/��"1_H�ʲfQA/���I�`卣�)�:��j�L�Ə���q.f�E��*�0A4NT�x�K7�|QO�w����[J���h�ɋ���3{y����S���$���� �@u�1�Fn� AmE /LE�X 7�����#s�"��ZG#{P�wGep��L��� à	q���MK���J��?ƈS�F&��6���s�/�7�[Hylc�Wl>m��#��ED01��n }F+a.o.�m4	(�u~M��Ҽ����2]nX#�N�%:pܨ�����1�<�����B���fD�Ij�,�<�e��@�
 ��i&���5VI��G[2o���&��L˒����h�B����B�`����A��ϫ�=��� o˙Z���D��f��$]�7���|�3�WˮuW�R�M�2&����{���_ �ҝ�+iD$L�2������]u#"Fʜ�Q�	���k�0d��d�VR�3I)\�sW���e����uPߢ�R`��~�a(b�6!�.�;_Mٓ0R9R��S���zfҳ�+I �a4;}Q3�AI���b�G�y�8�4�?�^��=�t�7F�����d5藽y�"+�J�e��2o�8����h�Z�
 �ڹ ����%�v>�	7�s)�y>YI�������_fs��Ot3fϥ���[d$֬ϩmR������!���R�)��ɭ��1�ㆌ2��F�3�!ׯ�e�����5BO�0��sZ�Oc����1�M��b��}��ά����P������V�9w2n��l-}��WX�l�SX��L�ƙ�u�u�J&RGyrsb���)���g�n?_V����Kܒa�I��&;���o~�^V2���ʬ���i �ט9w���#�I������P`p0�b��^�A���Ġ��A�ǌ!W���{)�aWʀ���4ŻK�Ğygǧd(jik�z��Tzskk��F����	�en��c�����R�7kz�����o��;k��k3j��^��O��m��p�q5����|$�e��J7����@)����ά�$�^�ڇ��+�Ge7�e6�:�'ī���(	#�s@���ՙ�n�Y��`�gj߄��i��P���oo��*�L���fZ�C�I��>��y�.�j�UW�YФD�BsK��hb$����~x6uQr){��G>(�<��>G|�2e]T�驘.b����H9|�E[O[�GT���
�dm�|P�4�.{_	of��fJ�U�*V�9�	PbM=���PQ0��02��#+e�q�\!����m_G����"�	�!���'#C#>P
����p���3E�&�LF\�����Xlԓe�p8t�k@�ԁ
���白W�^j%a=4���O�}��ٜ#�鉺<���&R�^)=�a��J�RY��}߻/qOĬu��7y�b-}J}'	��&�ap?
;9��sGh��	�Iۏ�<M�ò�X.�X	/��=�ӎ���z$P�8�&'MOsħ$�9]�J�dK(`[�?@�CI��`:i��*�@�gw�3A��G��IGŬ�hj��9l����
����`Rmk	A�qQp��mMf�� =��d++<�'M"׼LA��j'�6P���a��߽K�<O���1?��K���-Y��^�6��U��6�_$�l{ksv32�2��]Bg?�c��~���o�}�[�jN�I�OP��� ��GV�DQS��tu։���{�<E�>߬0nn�A�C�2���[���u{��<�tO���P_ǝC����#��㜒V�u��8�F��In�O3���簳�XtE$Z^㙂-�62	�Ey��)�Z��Vް(Y��)+)��R�W,��L\r�\�]k�at)n'>����ӱ�'�o4
�WyR��e6_�،��	�c�n0�Ml._�<�gR���Q,�RHvu`�M��S�/z�@�A����=�8�5վ��=sE�'�>�a>"�,ޱH��'���s�y����	C�Z��e�9�!v�NM,�P�����!ƻ�+�)7c�a���=��-���z�MK^�Wʻ����Ua�u�5�¢��ve�3w�8�W����酾w�2u���?t�X���0n�x�qz��Z��k� ��;/:�4�.��a���,����x?�R���z"���C�����
}4d>��떾���Ҕ�|q<�����2�JU�[�x:��oR�MGą�Ν�F��_�4���C��վm�6�޴�a�i�x��h�� ����1۶NU�'��@UT ��>?֛��&��i��~�b��;P	ӱ\�� ��o�c�L߮����U�8�[H��qD\��t̆��R�d��i�gh�~�O5�:>&�t�Ǎ�@9��4�"���NN�e
�2lۆ?�TN�f����k��m�N�@BQ�ǃ��8��gz<� 7k��.������e��� i�_��Qh�
߇:�P���>��4<�RǈW%0!�9:��`��=�ľ�������3�3�oy�E2�-E�����f�U�Y�����z�G0�0�Reԫ��{�\!���^���s�18
�����h�@����h��,�	3����G��= �x,/��㝅�5Qp�%df��KE,A����΁--Qَ?3Y)9?^��O��Qh}��2Ż`��P�WQa��-�a��V�y/L��Nx�?;\ӯ��gO
E>�Yn0K?~by�s�&V�����m7e�@��.�;��O�!=����p��OJ(����r�O�@�%Xȣ��-TH�mK����"�eyJm�֞����%_��"z <�@������^�_$g�ƾY��P��4˦LL�s�=4����4mң/d2I�0E��ދa:R+]��z�M�t�2=��7K޻ǿ� ���c:<���7����:;������,x$�v�nKT�z��T5��-"�PK   ��KU�р0G3 �	 /   images/c35f35e6-9335-45d8-b9d3-3c107d870976.png��TT]�6N) ����ҍt)]��]C%���t��5tà �ݡ� =�C~}���[�����w=�<sΞg�}�뾮{oWS�ŽGvW^�:

A

N�] �����
R��B�Sli�:�V��(��=�]TB��,�/
*ʝ��((Z���so���W4��u{E�m��-
�_y\P~��y���ϧ�������#

z�������r9���ǩ���F1E��v�����?���Z4����f��㮣�$T�nj�lf����O�"o��[GKwS�7�N �7�O~��o�9�����n/�DGY�F��͒�������=7+!�2�D�ظ��qpxyy�{�;�Ysp	

rprsps�9�@�N�o؜@t*�O=/,A�n�.��N4�Ϧf��O�����ϟ��m���%'�_�:�q�;'�?z�ϥޘ��)$���Dn�Ru��^���ĸD8����j�v�4uwv�tvv�������O�9��~�T��FU�P�?3$vm\�	EE����ԝ%lw��d ��{�%�^�F�(zy/�^��ڔ�3���8Z��>�����Q6�7�'��
7��5g�����H����B\�NK�N*著���*���~����a`�Ɣߙ�����R� �'X	����
�<�ŉ��/ay�`*�l١3����YT|�����A7�� ������pFY_��<��Q�\$.*��!�����b��V���	�]�hwOM�E���9�o!�|�hX4�(��嗆ɠ������P�k�2^�e���P�|�S�h��ҥ}_�NTw�<;K٦�{l,��k ��]��''��H���{���<��J�_q�Wea+�O�����x�%�0�"��e����"mý\�����̯���yn"x���{DX���l;�c����af�z��mj�N�V�1[��K��̂N>�:X��G���1�Ż��ޠ ���_r�{(�����'�Q!jY}�4�Q���?\pZ�<Nv?>N@Ak�"���aA�[�l�3ݿ9(hN؃)�W��Q����X�(�D��U
� ,�MΌ.w⊰��؈��Ȣc��"��l1�L&1��=`�����K��� �&	5��@��%v1g��3���>���3_Ͼ[��h���R�d��h|�)lM|`f���KB��4L����/,e�8U��-�̖�K��Ӑ�W_@"+����{��pu��z��i|�<I.��i���͚����F���KB�#����ن���'s5V4(>�g��c�9�WH�x�P��B���v�j{X	/iW��_F[l���W�%	��a�����C������wC3�)�)^�k��kD�-�)$�'�.�_�/|�����Iq;݋��+3�0s({5\������Z�u5��@1�W.Ձ�p�D�^}���b��C"��>�b¯	��y���w�C^�(�Q+Et:�9H<B����p���;Jh)��\7ߣL���w!��7ە�PO{RE��hmZX�T`Σ���|x���b;p�].�_�m�>�`��"�.�~���ir����P�w�("ƶ&M�H�]\�XeGD�#&��+���Iť� �0�f�^����zǼX�,���I����.l���`��#]dڥ���$V`ُZ�V7S8R��ͽf���[Ěe>��/�P<��OR0�z�*����j�=c�e����kBп�$�j��t�uO5C;�q2K4UxA�<���i�i/�s��R�!��'6�m .>���qY?����a�������[�����?=9rE\}c��&����b·>�+�g7zZC47�kʋ����37�8%�ݓ�6��Ѷ�XRf5SVa=C�4y@�?9Y��{�?y��T><0��V)=�0���w�c��I����iw9��儑uH ���ò�C�뽜�����fqڞ/��R%��$Mk�e����7���d6t�D(U�L9��^��<õ��"��2m������6V&�<6�S`���cǖ�5�S�մz���Y"1�d~~��<3y>����l.��+��k�.��@�@�P{�l���*��]؏��oؕSFNV�Su��d�3����UM�-�+������?$�=���j-��g�T��xSʅ���SZ�n?��@+��YU$Zl�K��*�\�{�ʷo���P���1&c����g��� 7�`��3��Ϧ��V[���i���";~�Q8=���V�� I�z�e�A97u���%�c������pEX�Xz<��-��"�5�����N�y=��()�M�}I�i|��]"[�f�c��6����$��.���
7�ܺ��"X������Q�%��7(���w=�Q����P���˹���Nh�d�s����[�y���8S�F���������4����o>uU��l3mLnR��Xmoα�����v�K��3N�H��)�X����VNa&��
]�+�'o6�?�O���oŘ�?�W�J�K�<D}k�Wp&�V��]��f�>BF�W�^��7��ybX=���a����^��n���p
����+��uSK`)���69ԈS^�.lTF�l�2�����b�4�[�ȴ�����_[��&E�UO��f?�$�7�[I"�OV
�zH#�6h�����qD������9v�ˬe��
ӆc��D*��Y�����!��D$��bţ��H7WO	7��?.������DV���������L��6!�PB��@�M"^����Pq�WY�Pf]Y�o�~3|M4��� Zz'�p_ؖYʲ��%+�!����{5Lz�l�N5���p�\"���ѻ��^�+'�� K^;]�~�y��zO�Z\��Y�k^��mQ�y�Z[g�%��ϷS��:��>\����i��r����b\�[��u�ݖ擢&��:@�9_���ɑ<�|T��g�	#�^�!r">��%�RB���Vp����t��S������N���?^ȃ*%����I=��G��$��=j�<ȵ�(Îs�w��*���5y�(Y"�E�]4 �1u�B�k�`"&�� Վ~M5 _tm{���.��J8�6*��z-.�:p��[���Ǻ�?/:�%��QC=�Ql=O3�pkD����m��5G�ýs�����x�'(e6���قn�p�F�u�z];��OsRދ<��
�6�W.�̼7&��7�<#@�D=@���Ʒ�e�FE��h��H��V�u�ud*?�0pY���p7�-�.��۞�L+H�8�Z�/���dAR�����阑
�>��rfO��L���������_O�g+8��1�v�"w�����z��{��O���d?ۏ}����wM�����ځ� OD��!�-��}�FH���$r�Y��t��.%�3'2b��"�h�(wI���R�4���%��t?@,d%����=O6Ģx��7穌��vF����7��J{�}�iB���U�A�[;��䌖M���'��מ���g�[���]�Mp TC�]5��>�Eߴ̝���{�ej�v��-�;�[{��l�쇭gF�yf��Ҝ1�i�2�F�?ʱ�HS�-u�{[��|!�\:5^���t�*�m^tՕ!n�P�2h�ii��U����as�<�9=�g?��lW�ߎ�R�(�b�#;>u򃢬�g���-> ^/�.X�8�A�l�}�+��N���Z֞�X�Ϳ�eNN��r��Ϧ�6���o{�7�ݺς��tvą�D�)�5�wΞ<ѹ��n��S:E���CPp�mK�7�]gs���j5���]켗����R􄃞�����x����;�����!Y�u��
������K/"��F�E�v�}늺�_ȵq΅�:;�z1!��K#n��V�t�F�;hІ�����11�1���oǢ���W6�{p^�=�7��#�b�.[�OM�:�R�<�o�i�G�Wx�gV�?Zm��L?1��у���B��lA�B�X�&�]v��{y?%�/1Hq��:Wp�-��#�ĸ��4�NFYs��ȴ��2����!l�A[۶�����a�y�
_�3����6��g7jV%�����{�?�hWj$-�l_��ߠ��þ�l+���w�ˍKw��q��L�M<��x�m�]æ�W�U��:��Č�q�^��f�@f�1mf����˶2�`R�E8&��i��`T��pф��5�������uJS��t3�H�r�˃��%틓,xb��x�)#���?E��OU�[��d�َMgQ�/�똃���|���l���KD;���/!�C��~1?dp��8��]�s�^�9���3�6��d̉�t=��tS�L1�vZm��	#�[P0p m v�m�QzDZ�聹�bmb�����&��_-R�A!�7궂�[��f�Z��+O�t��W~`A>�'8Uk��9�x>.��Y��h�&ȁ%�(LbԦ.У =����7I঍�S6���͸oe��>�Kv� AS�D|��/�B-m]A�=t�t���䍈Ր�-�C�&�Gy���S:#�V���!�ŀ��eߴ�e@����~t�a���j�7<A,?wDj����1��b����ѯ�)G�P&[ *��}bu��Lr�7�ֵ��i�5���oNd̡|�d&�w�f(�gG-sp\d�AT��/��=(�T�}A���f�i�g*$or{����l�(�����A�Δz�]gT����iB���gc����w�ϫ��e�e,�B�n�E��a�NԴ��N%���o�ى<�����Y�>M���'5trŧY�X;�#�9\m����+��ʊ��%�8U����J��gPl��HX|�80�t5h�W���6M��ϡӽ���!���,�8�E���yul�םt=��0�%�惏�KKd.�ٱ)h-�>7ne�2�|l�����&���w�!��7*?o�s�R�6R(��h>Y�6�l�+WV�M�e�+�<گRE��D���Z����q��n�i�9�ܿ�#�����>5"4g}��ug�g/���8?�b\G���X�E��[H`���]�:�k ]/Zѷ:\އ��MЯ(e^����n�^�T63*����1�/6b�>b��]�����k�xÈز��������٧�s�d��]ߔ�~��N@�5�V��I�A��H��l۲�5��D'�{���*����!�G�[UZ��=0br$r4p�A�1���!4J������F��b���^	�s�1)9q�ijSCc�u3y+��8�����	�y8���i7�Y���Ē�"�v #�d�V�]����3&�;Ъ�h�#K(�d�`�Hk��6yz�{�;��P�s���	I�W'����m�X�<�z"��}_o���>sU1���c�v�f%7��:�#\��Ure40Ӂ�E�O��p�0���^�O8$���)�i��.��L�ysJ�*�\���k�V
���bCR[��=.�N�G\J��)�xlZ�9L4��܄5�f����%�mU!h\N��;-��T&�7��l�K.|t���*�<�rfr�h̶1�oc�T��瑽�r �~��V]	�9t��!�����$����nh��>`��,A�[)��YVRc��2��nt���3^�J���ݐX�����r�[�U��l-�
lm�J�}=�?�4M5�3a�<m���xxVǗ:���Wr|f!vW�x��KL�Ӭ�kҐUe���]��	��E��K#s-��B�R�nm�WM�@�֖jD��̀81��hEd�E�5��엟%�<�G��{�O	��wܹ��I��t�Vk�xh󺲱8D���wkYηFç�晅��g�g#HG�	��GEh�ދk�Ї���n��xޒg�zƓʱ��^B_��l�*�!�`��L� ��͸/8*6�JP�;�x������vFe+x�'���*�>�+Y�?��E˶�Ѹ+�/�i��YMfض�x}~�>�.n�_��[Y�;�k���$��*eL
c�uu>N�`b$���z.�p\��\}e`�^Q�#d��DJΙPJo۶̜��WzWN~�?}�0�լ�<�H@W��'(�����G�_E)����o��Kg���%:m��^�h{��+��oP���0Qu"�$u��� 	�V�h��j� ϴ������xĊ_���~s �K_�gy��	ɨ�qOr�i�FXA������6�"Q�o�ߧ͏��ğ�8��*|�Z�P���{�~����ڶ����g����zW}i�0%ۊ��:N�cj���ߦ����D����������f�%>��Z����>� �`���C6#`5��+�AUwn��w����]�Nt�f�8<Y��^�v��*2G���J�;�x��u��A�o�E������2�x��)���]�b���}5���~$m�$�f���x߱�٨H�`��&p�M+%�+�r)��Q����\�7�@Z�'U��&;R��s�K�{��c�����v1���F��[�2�T%�8_���|��NN�^���T
��ƕZ�~��Z���6/���rԁ��<L/�����PE��&4Vl���y�UL��1���&|�3e")���Y�}�M�1�E;D(e׃̩ �-z��in�ǣ��̸Ñ�I��Ƈt�8XY��8z�c�q���W�I�r�P���B9�+_o}��Hp�Q�@������x{���޵�[;o��:���yͧ]�}�_�l��m�PK1<�v�{��F� ��<B�h-�h���$5��@�@�ɇ��i�Ua�x5�!b��'�k��g61Ʉ�;�㛲K'�<�N�a�l=#ě����~q�v���p��]_��'�,��`�|����F�I"���~t`�����)�+^�VX���63�%"4ߜ3Q��۟M����{�m5H�v��M]��~��/89���hK0"l{3 {;ɷj��,�`w�A�s<��p�1�3>�j����:t6t�ğ`.���3��5JxU���e�+��|�1���#o���n��xO\X��!�`���B��5V�<:��y�+�n����l:�i�N3����0���P�O�u����~#��v��%�R!��j2����0Q���h}�e�>#]i3����GN���}���j�ηY�E[�|�qҬ߇қ�o ]�.C�Om���\���	�{�|L���̨�f�|UO���o6�FE¹!;�r+scd�y��+�	''%f@(哸�L��x+{V���9������cT��G��~�K�PC�yG�675q��֏W�c<�{�f,s:a!�.��\��C.��|�ٿ/��}���zŁ��ŧ�J����{C{���v���	��-���1��cX^�狫�}�M�|'�b&�^JzY�mSj�����p��Pv�l�����޿V,�M^�"W�B�g����*	�[�O�þ֞1"��4
W�S-d�Y��Ӛ���}by�����^ ΛP��y���b�|�� rQ~lFh�=���?Uy�܌{�ѓ���~1B�8���r'P�m��'�M���~>�?�M�'�E���2'� �2��@�i�O�m'F��,`���+��	�@�ͫ��(��ub�c��eX�5��>�����[�+|�2FM����
6Z95����|�vV!��$7�'�hP��	������+��T�Yv�kz8�xu�k�R�!lg1�^x�(ac@��J0udL�d����ϭĶ]d�S*����֩�^46�ߎ(qb��55� <��˔K�Ԇ��]��Q�K���V����z����-;��k�(=f <l�0�n���)A:aݑ9�_[�k�d������;�*�j\�%�O�f �;<�r�l?f�v�9���M )���AIC�A�g5G�]q�Z#B�9�
wՕ�TaXSm�ʯ�g�H�e�������4�:z r�>�:��L�ki4��h+�J��'|�����v"�����s/��BlUU؂�_�;�GS0��_��Դy{�9����(K˒�}j*(XG�[+��W-0����-��l|\V�V�w�\Z��1��N�S&�8���7E�ʧ�b~{B�[�3�w��Z�A�6�fR+SB:�����x?�<�Q6f�R����%wq)_ݫ�d9��d¢���~���K�O��5��q�/9O���HSڌ`m<�9��Pw'�����G1!��l�#Rz/�H����l�x��	����O�e���EsM���j���2���c}���n<IOph�`��9�4!�.k���n��Z|�j�]�%%#��+��O͜��1��x�>/��<]v,�i�Yq�QK�C�&I�J݄Z���E�a��Z~��^��>iN�����z	cĳ�9	mО��!_���O-{��T�O���m�+A���6��ƹ ��HF��H�QlB���7�=d��W���$�X'�򗚖ͷP�ѾW�b���KH��Y�).�)H�`v��s�����o�>�c�����K[�	=e&��3Ȓ�8_@Ė@~1��{Q�!9$�x�&z��R8�on�`��I�D���e�C3�a� #�� ���
p���\�hBµ�g�������{�Bu�K�>� ,QY@�?� ��!�M~,��G��q��VELh�'���EB94���(*s��P�p[ �����O�ͤ�O�?��C����iӖo�W!=[�z�\z�s�T��(�@�?���Pq�V?�_v�//�ʗ�*�ug���<$�jSm�6�wI�-T�dRZ�Q� &ϻ��6��yu�� �5�o�p���5y��o������B��;��c���w�Qw�;��',HP��-���|�<�oB�FQ�������\:�Ǥ'(�R���M����GY��ٔ�t��u^LJez��A�l8%6����ɫQ6!0�C�JD:��u�;U�(F
� Y!���DdY��Wl�.H2�0�n��>�.�׾��OlnjV��$�d@���P�^�VIE�M����6�h�	�x�%)��2;+�"���>�V�م5L�L^���Q�P����		b��5��fD(O+��o�[�4^�j�<3�k�|�8=�>�x/-q���ژښ4�G"\%��������������+�~y��;��~�R�PQk����1�ם�穪#�Y��0%˻�u �Hh��o��:yJ�甍m�&���wM{�!�����'�X��*SN��#^w�4�yn#\��V�.F���G� �+���$�w���+�EE���Dhtn�E��4�N\����_j{Y���ck#�ʕRE�K���p�Ȅ�m_���s�e]�w���B7ѝ?/��4��x��+S�:,�	?�XG���-2����J��-��2֝��f�h�f����S���ێ
/��x������3�	;2�t	�eћ�Ɂ��ڈ����������dc�co�Yf��o�A^��},_�[�_�,�6�9+q�6�#+ �#5��vB�/�̅$�l��D��SF���l5�l"mVw/	�,��U�f[Ч�;��<>	W�b�	��/f9�1��N�i�a�(�`i��##�5ů)�;�����M?�a�"��]*�\J��Z`9~�ށ?�m�������LK��7*Fp�9 �F��}�2��5B��͞�β������i6%��s��㷴ji�f!�(������n?dp�j�8mOT���Ç@&h�!����L2��M�~%Kzr�xdɀp�ȽpAe��̫5�̴�Xt0�6F��M�&�U�~pQu��b$f!&pcpc02p˧%�6�� q� �=P;`�It�����E������.7o���W'P��&�1|P������;��$��KW� �LGv
>���K���N�v^�a3�=�Vܴh��I�Mڷ��9�|��ƚ6��6d�׷da�s�e\>��(+˫!��xJ��+�5�&nq�܁e]�!v��}*ɨ��
Ùb"v$R&pA~�KFm�B!���8��j��K��������e:�5���8%~����f����[�tV&�B�ݶ�.b,�y{P;��6%�ȇ�g�9�c7��\����5�'9ox�U�^3՛��!�X��'/����]��Kunm5��t[%���#=������[˲�@�؝o�������� D�^�OL�ѝ�<]���i"��.���G�)�o�ό�S=�s�w:��ׯ����[���p�X�S����,m�b:�7�Ƒ�A���sF��-mz`�����+ �����s(�χ�"��u�w_������N��b�O���U'jKTp,t/X�4�7c6�r[9�7���%wRK�X= �4� j�-�Y�!s`7�f�KL�@��7~�Y<!Z*���m���a}��)o�cm��ka�9�I��<��b���[jI[%%�A$�Gr��W2s�˃;��rC�Z���.ܵ��CYWl*ԥ��O7)��A�r��w��_��2�����gjI���u6�3yYn�͂��z�FK[̗#�.X/�=��"�e��n0�.#j�>��S3�J=�$��@�����%�kY��ƍ&7C��kנ���(E�y_k��{��:5Zٶ����4%z�xEOe�y��U\��9w�1k�S�l@7��K$�qhB������%��1pa%�@J��#�����,�']pu�9�"��]Web�O���B�pW�qg���vi����Ş�I
��=��Ҩ�"p�y-�H�_��ԥ��K����ZI�^��ʪ���<��9�H,ڥV�~�!nd�QI�G����]�\}��m��9����NU��X	�h'~���2#e,�?īK$��5XH��oݳ��%�e�6�
CR�ݗ���'E������3}�aQ��4ɂ�nׅE�(\l���'R�뼩"J�M[7Q3Y}�$�N[`_h�U�c�zGԨ���ŜO� ՞6y�oȴ:o�:�Z>�7��GC������C�3G�pϳ<!��bO�Q���owg&YC�ע�I4��~4x����~�XW[�3��Q�I� �|��g��d���芩�ߏ�G�)ǎ��o�5�o��$��k2�'��ˊ$Wv�.a�3Y��e2�'�19��e��O�\��K�"_�����F��G�
�F��?-P*\���O0�XI��N��BIo�(I*5���@B���5b�n��e��߇�I���͜-��r4�%����f�A8I=����P" C/���T�e��֬��L�S	�D�'��m�'�����]��3�Z�MM%�<0�/�+_l�mO7�� �nU�I����O!�܎��ݪX��i�q +�����>���ө�V�|ʙ
>��q�Hj���Qse|��T
ՠ�P�b]g�lb)�cu�b�^''���)~#�Nn�=����ozR��a��%�q�e%���m����uF�`�Uap�?��$H���oӜ����Lx�4��K	)c��ޡxQ�q"��^�Uj��f����b�?��^�]� ��Y0���Ӟ����҄L��334N���-0o��Wٔ+�=X x�ӟ�ɷ�xe����%
_���mc6����d2Ӝ�G^~��w&���jPf�y�F�{��]�ktj���df�?���:����U�٢�᳘����K��-�}���-��n��Q�U���4�S�/�!x^ξzLH �*$#�0G�q	���P;b��D�<�V��|����xn���3�t[��j���:,�n��i�m�V��n�\]���'E�š>pK�~���n@:�d��T6XX*����6A�F� (���a�&S
���)�)v֝f�_��6���;7ߪ��8M���X@����;ɾC� {-��t�����jv.D%����>tSK?zZ�8��V?RX M���n���'g)5��>:�e�*��ǚ���'�!6�8/-�Z���)�%�J�	�BO~�3S]&���-,���6X��흘H��?ռ��.K�1C�Tz��X��
�~�U<Ե�J�]�� z6UU�eVmB3�؀>��u��u҆N��x�.=lNL��Hj;*+���I���f�֯�P��(���,Z?�7�0<Q�#�Z�(?>��WgU�Xh�Rp�$3h:��vN,���CZ�y55d�Z�!�Q�K���a�p�:��G.\[� ����'��^o��L�S}A��(�L�0�d�5�%t���vFn����}�t~� .��>U'��������G����_�l�������	��X�� h=5�_��NDЋr�[�p#]�,����y^�2ޭ��71�m~���6�sa�5�N��[��;�|�ȩ�4�����O�$��x1�*dp���Ko8�Ra89��~.�T�/hPS������[��s2i;��ت|7�"}p�k8$6�D��p��� s�H|U�E�#}�B���-%̲���w�~����R+.�v(��쬱Z@��e�e(	�V�pc#*װ*�B��YX�������R�X�UUk�%�͒�?D�C� ɥ�#��Е����p<g�yx/o���&[oFS���D�6]r���d�R�?��Y�M�W�1�ʖ3�Kf#���L1Q1Z��~4$v�%�t�r�"OwZ�6莰#I���8,���9�HO�X@�N�l�^�x*�"�j��RRP���f���34����TCÄ��㼪��#�8ߎԩ����Q��~H��U��+��F����P^���f�#r)=$J�CK��K2�=+N��"��2SD��Vu���;�	!=�bv@�s\�L&"�
�֭��Y�ek^ٿ�����N�s�NjL����i�S.��[��Fj3"<>x�'���LDeKʰ�k���#߲�ˉ+��}�* �ekHf��J�����T�o�Dn2��|S_���Z�L����I5K`m5���L�q�^��f6PIm{�o�UB�'7��Z�b*�cٶ�~+�Iu�����\���Θ�X~����a[�&Z��ߛ8hH�"{�T+P���.�4_�1k���Ie��q�n<҇�T��s�v��Z	K�?����1�7329p���rߣ)-�N>�3o�)�4g3=� _	O�#%��ң���i��np��м}�;׃#IF�C(�]�!�!)�8�ܜ�X����P�OS|�!� �ab�z�)�i��O�L������<B4�Q����F����r]�������kզZ9�)���W��$�:Z�Mh��<�,�ec��#U��	k����@,�⹧�I� �4ֆ[�2�V��uet8η�Ƞ�D�D<]'�eno��-*��m��Bm�p�8XN��nD�,�<J�rm�(�x��Hn���NG��E�}�]�!�|��_�ܞԉ`H<��T���'ʂ�x���~?��*݀�?mP��a��zkX��]L=j5�M1Jpyi!�����QNX�&�ր��{��j-����X���5���pg��nd^����Y�+�1��vN6�6�n����.���\j�E�]�?'��,�M��R��<�X;�����*?���� sɁ_��߁/�TP�����]���\���>�d7~�����ׯ;�����q/Z��|0*=��%��F$z�	�;-�W�ߺ̂�9�Z:��,��'�'���&KU�=eմ�Ɂw��M�`���;̦V�� ���bRI�^�{�K/��*_N,I;�Xx�~�6�
�����:�B�9���Ӝ�dGV�<޲�h����j����¬K�vM�ӡ. ���|�6xA��N;��\���8��M�ٱ��R��M<va�!#����bдEnk���� ���w�f����N[�Ȯ��!!����֘�	FZ�����?^�G���0V.��}| �ft��,����Nɚ�w�FJ-c�:5�q��b���z��}�ޠR�7Ç���,������a�a11l��f(AK�S���$N�{{���5��/?�8nͷ��?p���t;�ui5�Y����z�=\� ��ۀ^[ڟE��睽|f�[Oa�<V0�����O�F;��
(� �.6�
�=G ~r�<�`�\�B���}�俹�����{�X�h�^���L�{i�(��O�~h��r������?��O��e��ڼ�|#�x`az�p�9|Mam�lay�☑;���_����Bt؋�2�g�vou���~� �1k�V��-�we��!3ɔ��ܓ���U?zp�-��`ۼ�i���lS�r�k��*���h���������bK���v�,�+S���9��D0�����jŃHJH	����'�m�)V��òԨv^�P⁈��C����d*��Q�Wt٢�/_\<��⩣�͔�U �l�S��Q�ƅ������_Dc\�����k��˛�_kN{��*����B�X{�F{y.r����*/��D��㒾��Y�J�:��g���{Z���a�7z�`���5���]���O�{�l􆆜����GKA����.,��q��� ��s��j��J��r!� !>�Ⱦ��z��_VyI
ދ�)ߙ��x&֛4Z��߽w$�,�(�h9.�v{5��-��v�ۖW�ٵ8�~%W*�9"U� ���o��![�Er�vz��29,S�RF2��g���*S�̽C�=���!.����(l�Cm�zf� ��Ơ���O�[!y�$��9��v���H®�.�&67	H��*Jt��$���xXC ��!M��|ɗ�>��`e��6$��8K����e}4��&Ͷ�m�cD��D������S:��N,����BbI�`s�?/�ɔZԪh@�M���W�P��"��� �$���ts蟯��K�t��=�eq�h�[TJ���w�8�bL�CoL�1�ҏ&9$4�.36�0nl_�Ħ���=~��@�郔�v��{�[m���µ8�1����|����ؒ�s��w�+��[��l��5��B�����FC[�YD�<���$[��^u1o���/���wº8c�qڬ(�-��#�(y���	�z0\��z����>o-7Qւ�Ddt�8{O,���óT�l�q0b��\�^��6#��s� 3B��1�sI�ohRɚ��cMN�����D�R��~�T �p-�u!�#U8�c���8v���G�,�-�5�A���W��5@��݋SkZ�i#�)ghG�sb�U�v{�Uwd%|���iQ�7��6����6H�;$�'���6�O���S�[�O(�&����Т�,F)���<���4�7$��u���[���� ��_�'�p�-��N�;ի�hjT�$&!�e��"�y~zV�8�$E�A2ٙ�'5�V�f��������Z��VN�r-6m��UߝO]�!�8�#OH���q%�3�!}#c-O?�� [�#R/?�6ܠ������G��՛�3�|��Gj���ˌL�������F?H���ۺ���@���U�G�IE⍉�%�������ơ ^�D}a��s�w9�hd��Z�B�b�T��3i���>m�A����>�����!��w������5/Ҕfj����bڠ������槽��M��ٻK�F����e\ID�d��m�d��3d&g��W!ls�T(��ϳ�z�����#�TUm�^@�q�|v]�����$|}�7�t�@mEq�]�Ý;�Ǿ���Tc ��P�C&�[Zb���ȣ��d���G`������1ߊKH�7����G+�HC����#��[pj��
�yvB�m����#��Of�wȼ���dR%�Y���k�99i�3��+?.o��Ĳ5R�.��w�.��;���J���Ǿc�E��'�Ou�t��@�1;��?�@w�9P�������3��h-�+}G�OoYC42W��m%:|%m'e��]�����H���Vpl� \R����g�;��HQ�8h���#�E�f���(� �2�c��Qr��U��w�?��(��3���
{,�_�f��F�	&��w�~�3�F.7�k�&Pַ��QBs����h`��-H��X8߼yN5�oߢѥ��p����)����5�*����D	�-��w�s�F�wψ��̹���a��UM�l��t?��[�IC��
b l{��B�tlظ=��	��lY�,d�zpI����+�G�U`@h�p���Ib�= r	:I��=zZ��k�^����ϕp��"�A��֖�]V�Y�#��J�97���Ju櫷k�nտ��mKW��/�G��0��b[cs[?"�p���K������`=�M)�/Q����HB��*lc$��'ۉ[�\q$�������B�oy%���Y����}D;�G�@��Z�u�ԫ
�F5K�L\���4������񥚟*����|�a*���6(������w�Sꢄ���8y~��jl��ׇ��ء��[��{JԱK��2�2}?�<���L\	�I�����Y7%�L�FS*�)u �?�կ�1	��ge�Ab/��W�̫K��Z���i�Pf4�xr�I���|!p��"M�-��w�\�+{-� �m;���P����S@�K?7Ĥ��g�U�M��H0�~�ЏG������ŭ�*3� -=��/��?xSz٢�a��0�v>IՍ���l$�&*y��])� ApD4��N��5�sʌ���|�X��s����׈E{�er_ݡ9� �r�s�SVOY@'�xT���ଣ�>mpT�s��}(��
2����w���x����W��uM��V�
�S�Ʋe��5[΀��3�=���4�:�mɀx��sU����D���2��Z�4�]#I�_#�|^v���J=�9�h�{=;�k&���+	8h>To,TY�L��q���)2��-<0'��Z���4~sr�����/�'��Ӭ�^����t�^���.װz�B�*�FL�c�O6>*�^��鹨���ݪ�|������\�}r*ёk�=�"zHķ�;���+�K����V͖�q_U���I���������}j�1U<憪�������D�-�2��M��١/�NO��p��Au-]��a$���@pww\���n�� 6������.�s��[oN����E�Zm��c��^����ǣw�g���QV*���>F�+�0(��ˁ|�[bw�C֍�Դ�;+���sAu��"�F�*�o�U~V�~�W�����=�V^1���r��XG�_�.Wb�dJ�������!��C��[m�9�96��u֪�H�V�7���&��χ��G�Q� ��.9��J�tK�D�eGUT������뎦���t���K��������\'N'���i������RK�6�`�����T=�W�����5�sj�jЅ�"hK��B	�	tY0���~%~�3m%l(��������ɲ7��rn>���e�h���YX��jta7|1q��mx���>;�:CU������ηN�C��K@s�����ٿ�㧿k�2��m��a*ޗ¤�i�;�>Ӂ��\h�X�1ܩ��=�^����W톻�:��Z��}��	 �;j�^�r0���4l��9H�����ūm�Nį��8�=��8hK�"�l��S*9� ���L�tu���%I��Oe<�����|��s�7��m�I�:��Z��x�F���pG�0"��Jxݟw��I���6s8?�����9���@M�;�NxIsp���U���k�N.j������)�^gEyRe�}��F�m���s.�^&��e�����6��j���O��t���s�9S�f��Ѓ�~�<Wa�&٭q	�}�f��N�Cީ���(œ�Z�X��L�\��x��] �{�n�Kg���t�L�nszw�yg��ϬZ�._Bn8yAβ@"���i&��-(YZ�g��'��T�ջ���3�~E�ǖ�]�M��2W���M<��g�d���^j{��bbWi����`���OPIyBb0˾&�,�=�:��G�
n7 e� y[0�V.���4��.��<�G<yfڨ3�:�7]ڃ��P��ʗx��b�bYU�����r[-W1kHS�>��p���T��-6Ғ�NiRɀҶj�!�~��SU3
%�ȿ�$Y"
X��)D�أH��mt���[�%�f��x5+/�� ӄ0�j9�d�͗�b�D��q*�t���q/�^�,��xy���E�/מ���^���������,5TFNċn�q�f���B8}N!�>W�n��(;͇���ʫ~�$i[�S-�X��):(=����Ţ�rq����F����^h����G6����G(G-'��hF�@*�h������C��a _�N�}�}�`�#$��顦���X�����)�U[R�)U1>��go�����غ�P~nB�ޭ%���"�3.�M�c�k*��Ic�� Od����k��`)k�� �GzJZs�hے�N��Ls:~��7�PkM1\d��=���Д��}�m�%��Pc^D��;�3�mJ����ދ:��}����J�LHq�A���������Y�<�>�8����oL��6=j��6��Zx��#�
bm���$�N���P���yQQ��<�%��"K��{���{闍[��GɈ��KO�J�rq��[/�J�NR4XBy,�`�L��̏��,��n�Q`�F�gF	ZIRP��6�ku_6��+p�~s����t������|Bo���H���L~Dk�x	t^W|� �Ф�]��7.���&0ܧ��v���'��m�U,�̧o�L"�H��B�B��b�8m�&���Bq�o�F�|�0⩯��F�~c�@޶`����S��9��6�Y�_(�8}��ӽ�v��+hkA�����|�.��	!pVc�VO�
�����T�����%�8���Ij}i�q�o�������
�����o=F"4'�w�U��sX0���?�Q�*(�d��pi�\U�׀��<�wH��'�bw'���OMc�r9Њ&�������)̿eb��رL��qC�NFV�D��or�Z�O���ph'Y-�sVg���#	LTӹ�x_Y�n#V J��ږ�{���� W�0IU�����i1��w^�k����[*A��N�R�(i%�X�t+���e��z~�%'n�zxY�( ���TF��g$�y�^����̣:?-���7��ξ�|�X1���_�_�v���~�; �k���Ȯg��ɽ�A(��"�讦{A!L��hWP������u�������E�b-E ��m�2���˾@.�OK�|A�(6�Z�i{�����Y�4��7���S@p��@4C[�@�3sT_X�1"	�13���,u���-31Km��>��5;[@�jp��p�u�z�8k�hV��x�ϸ��9\����x�p:>��C`{���L��Mc�p遃�VXo�ݗ� ��uT����?V	�Ejc>��R09!��eWi�<�̙�m0+az{�;�����l�08�Z'�?"�����?�����@\9��N�~��} �s|	��].s��`?�5��H��&�N�'�7�UD%|��1[8ٟ��X���i%��g-K�L�G:u�T��Yq�9�~d�?�4��y��������3�u7&�M�5h!N������
g�N `	dL�Z9z_�3���!x\%L-&#a-���8>��տc�ř��&IAϼ�ub߃��dҎ>~I�?��n��u�{g�ݪ:���f=��l^a�%�����Sq�_�?u?�GE �Od��&vk^X��Qry�_\D��r\�r3�Y�*2@b���y�������=:�*h��bM[e�'ٴ�O�B�&8�9���|T[�Fjq�7�Udx�Ä.�D=F6NBy+¾w|pL��(���(*����^�͔��G�X�{|L �ch|�ަ�V8'����X3�̢��Sl�����y�����+�̎��a��Wۧ82���K������X�9�vV	0�(Ai���mU�~?8�[��2R��nߪ�m_�o�L�z�������pvp�Ʀ�$�����g�m�t�ੌ�w����- tTKb[[*�aj����	j��n��!�x?�+��q��e�o���u/�"'���1��XDe�x�;�Z�f\�L5ҍ�w�_g��ޓ��$|$����hB,��w���w���� Yd摱/O1r�!�w}�Io��*�Z-�=/����%�-��].ʇ8�$��S����oB���c�H�.��"��Y�%m?�B-`���ٛ���B\m��7��X�Ͽ;Ӷ\�8ߵ�`'}��"u%��M�ާg��	�[�'8�9��T��Y]ZD��f�æ�?�"T+��.[7n��̪;���l�qL��?7'�ol�US�'d.�T��Ƞ�7#�	r�yY쏖��/.aj1�!4���w��`�����/�-����k���e������̘�Fux�]�T�[�\�O����+L�;���q^��O�Ң��Q<��/�3���Ϫ<.��f��G�,z��]^+!���6��{�4����	��Ȼ`?p�3�,�O�|	�s�_��PR���S��- �b��{�`R�'ԙmd�$� ���yӅ ��zs��g��{K�ר�N�U�x<K�������ǔa�B�|/;�,����7��y��T�󦒶��ޔ����, p�Z�>{(zҡ�ˇd����q�O��5��K�������n8��{tW-����տH"�[���z����?�,��s\��zy�g��Y�+��J��dgRNjKagk�	ࣕu�b�<�Nx �ߡ�~�,��M�?����'���9"�s��m��ߠ#a�/(�4��w��s^$<����iF�HA�����L+���y O�8��0{tV��Ű�y���ol�v���� ˅e`r�o�$��i7��F3���0���T�d��W�Z_�h���Hr��(J~=S�[ -E���s6�M~q��.4>���ll,i���i�ܮ����8uqe�Ñ]�h�/��#_��Rc�a���VECS�]�������G+�M�i��6�R��93}���Z�ї'�;y���x(��`2�r��Ha�"H{h~��N#1q�nʶ��o>pi2p?�4.e�+Y��.B�#����:-.Nu𒲌������~F��}��S�L�6<�\�֒R��#����WR[�^$W�B/� ��f����ǽ��g�����n�ǉ멛'0���2�B�nZ:����z܋쓈�ض�;hq��P=�Η74P9 7x����#�q+�@>����&�Di����z���UW���k�!$��V=IO���~9����6@�����P�[Н}�l:��)���7+��V�t�����!|0w�HAu�%Cw5?�߸L$�-»(��=�V�K���G.6�ð��=XMV�
g�,�z\���ͽP;�7�8*OS��Q��4ò�4o���z�$��D��%�/�����޸k�N�Q����,�=�ܬ�՝��3ʙ�߇�&f2���<�:,�`_�����,HYōmm�'dW��6Ȓ�u���ˍ��f�\��AAK�1u�h.&|!W��TI��f��A)���mx�`ymU�E�W�?�{�ޟ"uu�G'��z�qt�T��!��8ٚ�՞��2���ߝ��u�5]n��Id	��rJ��k
���2L}�L:\�Dn�y!a2I�MK`�����[�2�A���|Ԩ���Q'ˁZF��z.s��ۤ|�W�u���?�ݕ��l�eQ��B	�%κ�q��VgR\�͓����YS5���d�뾅9m�S�UE��6�W_hmm� {�@�8^�S�O�~�$�����٥]"�I��%*Rկ	��+�@ц{�Ӂ�(�F.�o��3>K���>���qXWoO'BJm`�P����Qo�&V��^pqr�9�ѠM��*��(_���Xo��k[e�qI�~��֝}о�^z��� es���^�w9��kg�s��3=�'~z���?�K�;��O�$�D+pa���4���[�^z�iet�F����x��QI�`��
r��2�N��I�8-�%��;~����v�oh�θ��PhPl��B���FX�׺�����h&}���7�/gR��=�ٴ�~o�Ø��b�Ut W��nwK�7E�i$��u�'ŝJ<��%�R����k�w簓=�!� e9ԁr�����6��$r��6����"���zZ[�_ߝ��򘛘�`�;�K�d�H,)��fƔ���x���	�`�ͥ:�V��'�&�������&:��W��j2r��L��?���.���N2x4�����,PGmV��ivQ6f��66�����omU�g�Y�+�AT���g*v�:_��=�%~�NI��W4��� .�[´�TÚkޅe_�n��R�r�45p�_�}�nX�����[d�Ek�VS�S[��o�?��(�=�*$�K�a�\V�������wǤ:��=��52x���	bX�Cfr�H}�Lj�e���l�"Վ��	nV����Pc��J�*j]=龊���
�6�a�5� �ǅN�-�'��*s��AϖK 6�W���l���;�:]�!��/�!U�J[���x4'�iY[���w[�<f��]�'bx��_�RbkHU�,b������އQxy��z�͒���t?����k��l�Z�K����ݮA�?�=���Gqm�Oh��i׽k�*߹3����s�`s�UrVz�j��	������I`���(���u�A�z$����C���a�rR�f�u�7â�װfkr�1/hVe�����Z_��w*$��e
,�Wn�M����5��^�S�6~�$I,l����r\�y|�<6��lM*�XT��6�vC��';\hȳ�Y����hu��7I���$���	�x��"����KY�Ŗ3���_[-k2�vQO���� >�x��zBn��]U��xr��RկxF$NtD���~vՖ'd�J���XS��3[����T����0t����/�faA�G��γ��[�q�X/f�b��.��?��;�IG/F��6�sj��[BC}id����Y�R0]Ģư#m�HO5�_�8�.��;��(��님_�������������ů]�#p�5L��_��˪(�k�Y���QPt-.�:�]ES��[�ץ1ؘ�w����9f�#!�� ���P'�P�2[;��w@�5LΠw<����k�h�X/9��ٻy���l<N�?_ �}3C{���*;j�����>oo��ҍm%^��|�u҆3Cx2!&{�g�QO�͒�Hb���R�]�)G�P��=]���N!����W����	���T�b���8�ߎƳ���7u�w_��jऑ�wpN�1֯�O�=���(�����ť�p�5��Z��Y6�T�0�r�.���1M���{w>��g�~�_��v��'�1`��+���+I����$���9�������.��p��*it�����h���Jj����sWђ�D;p����b�k�����/ǭ��zN�ݱj�|Bl�[n�iS`������%�L��4��lm��KK�#E�݌�z�
pӛ��I�1�F$h͉Y?�h7#JխI��*\VҌ�;>���A��3����8Y����3�q���B
\�����)�S��V����x�%�蚲:p2J!ޯ��@�_&ؓN��٥�X����@����p6��+��K�ؖ���i�܆/�u�I2E�5������)ј��YV�XZW���Jg����FY������Ŕ'�b�kwlL�5;�ћڻ=n�x8黤D��E�x���f˧��ᴹ)�\��0ӝ��hWqFXԎ�q���R��?��4,���`�^��C�d����w�2 N��Y������A*lȻ�Vy{�f*�i�J�)��1��C2v��ᏵS�з���҈�o�HY��͆��b+)hг�--Jh�w�|�20$�s�
�N&�1N{�-Y�9�96,`n�M���r�#��E�$�K��xH��y��6��~e��WҢZ�ӂ�'���P��o�pZ��Z/� ӳCo�?`�RtECV.S����P��&G�
�6k��j�wN(�=��I\/�"�^�cv��j3��m�0-|`|!"B۳��}�� ��SS,�v(�]��)��I<RB�I��wD��8=�j@�Q��Y����Jg�"�J=h�?�(82�vf�n�t�1MA��q�Wl��y��!t4�\�v�����G�����b�OM��5��8����"�pS�!�� ���z]��8���BX6ӏ\s��7�Yr�<��V����<�?�@�F�b�:�}�W�!�Q9�<���Tl"�q6WҀyN����h3d�8�P����@
|�V���mՆʂ��y����g��t�}�{A�-O@>���5("��#Ьٍ9p�`��_74�U�����L�̀\&@���������S��W�����-�|eEt��6�Q���_Y�֜���s�߀�E��3�H%�c}����<A�áN��#E�M�ي����E�����7$�e�Б�r�8@��=%��柌Dvz�&��jn��Y�Lɲ���GU�pn�-<xW�o���ݸ�?�!�&�d����N�t������=�����`%�����K����S\�?�I��b�{�-�P�O?�>����"Œ\HD2���l�$L�A�J+W�g�c�q�HE�h���3O۟��BC�};j����)����4���&S�Y,p&p��+uufv�k�����#p+��UBqX��:lk��^��rO����6i���2�i��gE����i'"���9B��)�S8E�I ��e�C�v�w�I��t��H̭�\�S�0���ʯr���}3���@v8��F<l���m�/��V2�ąt{&�E�|���lOۄ�h^W߂u���Q�G�� �'wFo7 9�S,���åbt{�b�<�5��}A���/a��u;�X(��|;k�2o��<G�Uz��=�/��^���oP��`@�r8QIF�^��d�{6�������Q�{g������W�6n� }u���2���v=^?��W+��ns����VX�p���U�Q��v{���ۃ�+7զN�_�x/|��^\$�`(I�@�E+WXYJ�26��e�����HQ+�H���Uov:銧[�w��6��!��:4�E������Z&�� �;�ћ2R�j-Ǝ�Bl�a��Z��#�We�~G��~σ�@�I1��5���
·)�9-�y�vڣ�`j �k���XX���8#-,v�.�U���OI3���2γ��r\,���c�h[���3SS4��\#jр`�Ň؜��氃`��K 8�F
ND|�VI_}lX���G����9�����	�;�Y�`e�l������!+"��<���p�^ʻ�< 8
����g�v�Mc�P���} �g��?�����+:P����j�>sSU�lo�C�
�0��;d!�$~'=�z�NjE|O�Ѐ�g������xH�Ru��1��V}��9�ο�CMf.��8j�b��n��Ei��4r�����SW�?,���+��)k�}��m��&��b�G7�m��J��+�e_������}�s��0_¸�M
C�͆��a�N�r=zO������3OM���̱�M�i�����ֆ"���/h��!��Hs��B��sv���:z]��P�Λ�k� T����Jѿi�D==�������9/�
�����U�iE��H����gH��Y�E�%��V���>�ؒ�"���A��"{�ul�M/��&l�@�Ps��+&kq�n�[*
�D���ɒ�/feo� ��-��&�Uݔ�m7`�S*�e��iӆ���&ՠh���hg�47V$CCQ>/~F$�1
Z��G�aG�sc��`����YIji:�?�Z��ʲ�M�F�pL�~���/V���>��~I�H�?xN��[�gŖ7G���@I���� �X+k@�R8�e(m[X\| ~��R1�͐��!�ϊ�|v/Rnfh�
*H��x�N� �]ߢ��i+2�0�?��
�!�E�$��^���}�����T��@F��w����cV�E$!�;N<{i�L.D�fֹ~��)��dU�n}~C�'��������sr�(��s����ٝ�UR뤲�p�_ 9� ���e��QQQ�O 9}����|�����[��{	�e�=d����؁��I~��͐�����ox�PZU\\�f�2���+䆵���=��v�9�k� -j�HA�s�3z勒��E�^277���C���)�����ki�ai8t'��� ��{���^�	SD��+���/�d�*������7��@/���Ht���6��-�j�c�~V+2Q��Ou G�kl�T2	\�{	�Րo�����鹓vA��WR�[�~�-OP:|���v�q�j׫ko�o�������;��N���He
�����a��`W�}���*p����}������@E" ��2�n�=4E�0���M�3�Ǘژ�H���`�Ւ��Y�u��O�~C(�"�RuE)���}�)����q�k�:��<�~X�$!ESK]����=����a�G}L����c���
HL	���|r��K����r���]c��}U>��U���ﴐ��jTFJ�R�� [g�* ��+��|ƅ5��s��@�t��������bHX�R]�=���z+\�2������}��o]�����$J�Wz�ls�,�)�F�*��"��j�S�9�k��x_�3�I���(�3���<��Xk�wZ�*�0�:q�0�b
 ��s��;N"�%J�?~8�k" LW-C�����z ��Դ� �%�2��9�|P�q1��h]*9����h�z6�_(��QUy�3pH����jqb�ƺ 
�Rkb��]�z��H�vK�l��s?���{gb�`�������!`襌ʘK�╇�����c�!�����G���$,S9������K(��~v}��Q��w$2�.'�O�,Lr�E�_�����H��C�k�hֈ���7�+v#t�[��gP&�o�݅sɯ��.���SD��D��m�mș|����!��?�1�.�9�6���o��y���d�[��Q�~������j-k�GP�)35Fk�8���k�Ջ�ܜ/e�����|��;��� ވr��Y�7�R��,�ۀ���/Z������E�r>�;k��h��o�y��-)6�.����F>�"$�������>�yâ��m8D��E.�DJ/�n1@�)���2CȚ:����p��q~y���_|�p����sղ�OX����I���*�k��ع������9�Hc�տb�:�g/��SE��7�a�|c<��vL�����T�_�xR�����/S~�f&@ �� xG�KQ�@�-#,w��{�%�b���>�!�3�M��Լ��I���U#�ļ����+���kRA޼����{G��/�S�Q��+6h�.��J��|��N;�!��݀����~���	�Y�\`=E_Lg�v+;��nI]�������ꜳ����t���$/�W\R�PY{	�C�R���l�V������
�m�ƇF�9����v}>)skG�p�YeI�$0�  F�>/Z�1J�׻�@3R$����:��6S+�U/|�!�tP�����ޙ;�ϲ���YVrb��5��ؖ1G�RQ��Bۢ�&���d��,�q��5�T#f�p�;go������)��9���ooVaX4�*A�wZ�?��D˺��4�2(=F�>��Nݯe����Y�Ʌ�|!qi�n�X��E��s��G�u�����K-���Ҽ�@jX���?{k��!�����a�	P�Ö<����(g|U���򪌄a�F���ͻ2�D������k)4=�go�V����Z�m�?�_��y�.(A�'�`�)Z�Ml}oÝ���!⿭rB>g�0jY�BJ��+���.��A��}6���Y�%��ᝰ[ʽ(�6u3����*��JQp���o�W�7�ӑy	�!l���$�æ��Pp�e��q�:��R��4\�U��y�ܜoU*�+'�Yw�a`�Ľ���>)���������?R���D[,` l���Wu����s�CX7��'�\���A��ϔ	�54��Y4�{7z�T`/w9h��E�￡�@�v��C=� �O�5Q�!�Re�i:e����q�Q.b� U�gȞǫä���D|jO�����8&�i���E(�a��*�n��:)�r�����4 teeX��G��}��Nb0���nꄖ�����n�F���
�����H��������K�_A�� �.���}o�D�Ż��W��g ��w��
x�x�]�|_i@}������w�?#�Y|��6W�uN
��6�=�o�h�2��+ۥ�S�p:�KP���{���"�VO4WҒ�(V�
nu���H��<P�6����*��N�9F2w!e��0�j���.Ru�+W�kem�Y�]�8�e`�I@5E������;&�R�vY���\��	�!�Q������2��g�L࠮=�������T�H�@��y��&VwK��"�/"����4�L>.꿇Q-��<��c����k���-�E6Q���b}hn���Z�K��L$�7a�}GEK|����������0f
Ʀ�zu�������#>�j�c�&(�XD �̓S��Q]A�r�w��zo_$XcM��_�!Bo_�N^�de��E���F���h+�_������iAR	Fv��6U+�S���}#�fJC�����G�>��Qo��+:��5�Q��Ԫ�t��`֔�
�}�\uO]�a�&n��B�i\�;��O��l���H���m��ʵ;6�N˟>|U�e����d��J��I�B%�QR(�+UWK!]��p��E�G�@|���������6:B>N>���2`A0����l"RǦfA">C�&=';'���ɣ���hV�����ܼ�>�;m�K�̝�-;=��2�Oni��T�F�/�r��9�z�{�wS0?�����؃-�+�.y������~�̐f`f^1��j�9��l|�HHL��2�7L�g%�A�V��@����
����1�5�;eci_�.>x��Iv�6��a�����g?��N̯{r�e۸	|q0t3��ۻ�-~�B:߬���[ݫ���b\-UjS�S�H�cG4|*�T��qWov�����+��!��2f�㕕
�5:�zs��L�C�∹=���m޿�'�%p�q�}��`�f�泥����/������2=
$�t��/�?|��p�ϻ\@�_�.�;�\;M��I	�:]x�mT����K�̳/,��*���EY��!�[_��z�����ƛ��F�Bp�k�ߪRo�c�0~����Y��x�nMMo�n��P(��f��q�6������-�k�i?��/&v=N?��Z��q~��l�;�pRύ����WIHD���pi�:g��U�}��Z�K݉��26�yj�4�= k����8g*P��J:H��`�q�EƢG����&����/z�� �_&\��h(G0��NS����m�W��I��1>ͳ��.)-!%�77�I씾f�,ZQ��<Ku�\���![x�7A?�.��^�hU�����������n��Pg�)^���(���u�˥�@�O�Je(�zܭ��2���^��O��dy����\�l�`F���LP��p7IǶwO��}��P~y`s6��;���c��IǺ��S�ǆB��f\ג�Tt������u�DJ�*�$�l�r3v��9,*�sȞhk��z+���������� N�R��ͱá����AU�gM����WUz:L�@�@�n�2��	f=�8�*rԄ����P����\�γU�^^M���F��G�-����m�(@��!/�mdJn��d2'�~N<��muFMo����#�:��*���@
���	�f_q�~X�����3ե�@�r.,"��H����k�ĺ15vX��"������D���"�RO!�k3G�g;��e�AO�Zcks�ӮLŠ�{ש�N��[���������.bZJ��ɚ�V����Ld�w�{{��Q^X�ч"���x�tGM���^���pYa�ͷ�ޜ��)Ŗ���G�	�X[k�錎�E��΅��~}��06���z
�y̎ɓ�~��ch"���<N�HP~��/Y�c�R`�����H/ūI�l�{|�fڌy�c�@�������Ф&��.�n
�N�z����p�w7
�)���_��>�񉻤����z�)�6�f�"�`֢��B/� `hi��3{�ϩT�o�r���AM3C/�t�2������fJ�ť�
��k�:+�O��89c��^���]w��ci)��L�2:�XC	��w<��ܚ�j�T���O�E�9���QVa�.�rh����*\�]'�y�=�VQ�-t�`�T��|񰕸c!�e�(G�p�7�0&B��BL��^l���aLR��ӹA_�h`16ԓݖW�/R���ɧ�}���I�hq=Է?��j��H���.��w��D��$��?����.�(�ptu�vDAxi��蘢��p�\���!P$�n�I��@19�BF�	C};vNP���*x��qι1�D��?�/��V�~��o7ڍ�0�AI1�'s|����ށ�E)̯C��(8;�7���v`����X��鄌�b�N���1�{�:	�P*j�O��e����0	��-�B��d�:����8O�����z�KT|�P���F�Alv���z��1n|Z�+EWaiŧBe\���� :��^�nzS%��:�(�SIS�L��N��W��D�`M��}�0�Ťf�ߍX��8m,�8(��~z����+�9 (��b�h.��e��9WTI�������u���R��;����,S	j�fR�p�q����ɛ���[��nXbxN���Er[��;;ܘ���6���0,�󼥌�b@}$��\G���Z�Lӓ{�	���[~�;�+1�P���եIV~/S ��!O���^5�Uop>g�0ބ��E�q_0����U��`IF��╀��R�3	�M�a�/��Ѣx�Jzy��8C�B]{Z�g7En��<`H0`HuQ״�2�UC~��#��u�;�:�QO�����V�]Y�IH*R��B�`q�g'?����o�9M�Q���8/s�u�,�s:I��U�l_� �/Z��h|�L���A�s�&&��Ȟ��kOſ��T�h%�m Ǌ�E��-<Z
�A�H�����n�{{J�]��5��c9aL�;��\ k�ͲP�_Њ����gCQ��U��s���T�_�&�`�A�b �k�ܪjG.�G�4�f�L�ր�x� w�Q����f]�b������m�oGʎr��\�F��^�a��[e!��j)��:�&���c!!Ҙ\Qu���v_�wp����Q�uD�C���w�c_�i#�4G��Y�Gj3�G��z�z��KN��T� 
z@�|(�L��#��u�&!��ҽ�Hm(�#����Kk�ƽ�9�SQ�D/�D%��N��r3`��.V�'�oN���wk߾6�skn�x�5��� �n�˘?�>"�I,����#[q䡹��n�a�<%S����85���V�+
kCX���������g���j���G�5FS���s�E�d�S�kB��jJLJ���>�^��`:���TL�S8{s�5�[t���|vϕ��z�V*b�:��P_��,���:c6 ~KJ⦤�F��}���҅�Iu�`f ����E���6�z���R5D�G?�fw�ف���n*��U��ܱtV:�Hm*�Q}�ʑE�����"x ��IYj����$�C�p���O�*���Cޯ8?����F=�Raa���`�����Ȫ�]�9���*<�.�}ť1`�.^֣��:p~H�{�j��V�f��i�Ȱ�T	�^I��d��Wn�\MB�:�����m  ����;�'��W����]�k�զ�j
��/�C669Er~)m��ƅ�Blѥ퐆\'u�<��)��yZ�p��F�X���!��B�m�:\�>��ѹm>�ʸ���ޚ��` �ԉ1@ Y�l�j`�̳�v��D�R+�{��Vp�Ӡ��ؽ�w}7fz [��aq�静���g����`���`b�����J��򸴱�������Jn%�w�-	%�l?B�_��n+�qwo�S���¡n�R����bXt'��!�Y�o��}]V�[ �%H�9vR��b�PSc��l!4�a��.�M��đS�s��Eː���p>)�k���9Հh9@�K�ꐸ\�D��@�TǰH�?�,};xb3W����- �5�}�l���R-)ߴ	�~�|H=!\ʚy%|����Qm�4�����C��q�L������.�n�����y:�g��L�?�K����GH�]��W�ޝ N�S��=�l]̏unn%�	�$�Yaۨ��\L ���E�_�6���2�h3���؈�<�v_�x;LA���Pr�,�饿�$iY�MBBJ�z7�|'Oc:/ 'ZJ����
��ȶ�����Hw���3a���"��wc��.��tf��� �j���2��F���!��N��U���y, |�6+��+��d4^�]fԛ����Q$=�硖**�a_��=4欂�� Y<�U}��N�B�Xo����b��P�?~�G3݉�X:W��A�X�ʅ���~��9���_����w�aL8����uC�[_x��ȢG[wOw&���L�t\�X��pW`��9BO�=C(�ӾVvsO�I+��������P]���5W�9o�ݧ�����j76�<Mx�mPC����[�`���mqhy�8N��v���ׅc.w�w�pbħԞ�o*�:LV� 5@��}����b�����]�F)�w�r��W�J\W��l�����>Q�-�Xt�����iu}%�%�x�il��q���ҷ_P�C0�x7�zH�LJ��Q���I���)�J�]�m��#
z�b���
�t�u�?��!���SO��<��ȵTwY�vp��US�w��9x4�����������9�K�R��زCt�M���� #���Xq�����������
����F��j/�fI�s9���)'�@�@|��'1X������i?��7c��u|�Qb?ђ$i���UP]ҏ�Sg&�@`�s!,��ԥa�<��ٌ6�+B�[�e(o�o�
��f��E8�z���1�嚪�K��D���.�Xtt����ĥwOo?MFS�{�~ZzS˔c���vṟ�)�;�,�;��Ͱa����z�M�b��r��K4P���8���E�ɳ1��1�o�}еD���Р*=ھj��݊v�{_���\��;���BO���g�}@�3�3�xX'!D�|�+h�I�ׇ~`Y�R"O�/L��ı.N�*����|�!h���9OeF}-&�tf���Ntv,��i�o�����cx����|=�!F���2��K�]�^��eB�/��=�_���k�-��>�3p�9�}�;�c
�ku�4I(�����c�0 �q�ȭ����L��C!�畻:�oW�0ec�6ڇ�T�����/r�Ls�=�HbS��4�Rr��5��0�H����]+n�D��Y��I�F,�[E�^Y�u>�����[8�������*-	Z�X����ol�.@�: a�X���r�!&k]� �6�-B���`I�C#v�i��w�9�c0��[� �*�JK�u�V���cĤ��I���������!_ؐu��wd����CG�!�j���G�f|p�@�����2�_�C��b㦜�$%���6i2ڐ�g?�r�|�e��1�A\=�rm���up_�A|	F���?kY�IY�go粴�L��!8��4� �	w� !��܂kpww���>��3���s����|�Y<�Ǭ龻��꺪��[���K�5x]���p#��O2�}�}��2�(\%m�*#��s�V���!׫_����d�|��	�ocs����ܜ	�
�1.�2ԄoҐ�c�
��$&U�f�E�q*ϫ{6�3/����鑱���-�D�_�����BC%\Tj`�����
~�MM+�3�eg�vb��pކI��ā�*}m_U�%o='C��X>I����Ys�J-x�"����[��&��u�?%W��g��[��aU�� �Ф:l�,�Y:Da�B�=Jb��9������f���4��t$��ܿ�t ���[5I��?y��NZ?{y9%�^���զ����l$�E������Rr�����}�R���9����a���F��C�-GH�m�"֢x�؀G))Z=W869�f�ڼZ����U]����"��)��p�6���8�e߻E�*�u!\@��I1<O��!��z�{��{����ۂ�6nIWM��bl8�}IQ�8,�)2�O,ֈ��&�s��P��Ɗp��ײ��v��h�$(Â�lm���B��J�w>�4���t��E�`� ���G��3,ȟ4�����UK�!�z�H'�#�&^$/��`-\/����a�U���Q_9%����?l���/���4��1+*z�X�v�>��K�;x����ǭ�#�p5Ot���o|+��D�.�������ғ�Yݯ�j������Y	��ʵ���к���i��î����=+o�k4���};*%C�%h�t"J�0ؿ�NIZ@/��BƲ�F���,6X-D�{�OuD�����~{R'q���S��o���9J�㢩�w��*}P��쎅I�liI~D�Ig2WY����X����zW�hwl�!�+zޯ�=%�oCV�_<�����vH`��疬I]��}#B�ܺ
x���T���h��cZz��0�v�K�S`�T�_d8$�a�|�W�E{�|�?D&�������y��X�������)�d1)��|Y=.��(a 2�3�nkA�d.H�a� �wT��^�Xz�������u�FO*"M�SmӝY��mdX�b�v�C�ªq��V��s�o/�t��FHxOF�R���]\�x���v�|�Uy���~g���9�L����z�8��N�N-�Z�:V�ة݀�f�"L�+ނU=�8����_H]Lմ�̊+�nE{�Ed�)���CE)QEG��y�-q��vH�h�V8��Ɔ"~����fG���U�l�1��{Um�z�9��L���F���-ʹ}�v�c��.����7 />nn����Ԇ?�sy���8F��<��7�;XB��8� ���9k�/*�]-���3�(r*=�"��o���Ϟ��y�L������h.S\�4��������%e�����K��V�D9��ВPPS��~�֫Z�ԛ�k�u+߁Mc�����*��e���5��GBHr9+kh<���u�\�f���$K��[Nmg�l��v��o�ԓ�Z����tRD�)S�*��o@�d1߇8/����]�j�bA��0/��a�;,��|fm3qB�����+4T�"�#��ϕ��ii�-I���HEOѹcCX^a�q�}��s��!aTvo���ޏ���:4&��T���m��p�S �,GM�TJ���K��ahh�l[��~���"�@��?A��4_!Qa�����K)S��X�ܥo	���D5)p��8���n�+ƀ��*d@�����j����o�O �Щ��Hb�w���Ӆ3��%5f��ᜀ����{!F�n���[hg4cfr���#���7���-撷b�馜��;<]7j<�+�m�W�.k�����e���p_�������:�>���CKsK1?۱�܇!=a|q"�A�v�,�eh���b�
�����������J��@j�#�/�E"���D��G���U�'���ݱ'ՋI�]%KB"��>f<ս'<�l_��x3Y�Of�JPNj'�
�A��!51���5�[�M�n�>��d�а��썯�M�L�p�^�$�&��(%oӇ�����2�-����9k\��s���*���<�P� �� ��R}����eH]�,~�3!^$v��E�~lG�fuC��fT�Yj�2Yl�&Z��Z�M�~|���Q�*��뼘�QY��ṱK��
3$�[a���%-Yo6$m�'�w��4k�?���m6��N�S��1�T<>I��R}ǧ�rf�(�8��g�j��rK�a�|$XJ�t1���*�MH��C���<�n�l�&ybn��=U�\�N�y��-���DS+:ˊ|�e'��9�n�۲Uǽ�K����Y|<GZ��U�{��b���N��6�<�#ù'��R��ZW�Eu%�֒�p3;0����~RM��D��p����&�)�4c��N�u�t�1i�a����\��В�8�H�E����.���tXR�b�O+�k� uwZ
V��)1݇��� ��ןi�q�	����L2��N�^��A����J1(ޱ�e7�zQ��>Hs�{�;.�+I���bYU�����|a.1�smj�d��2W�1T�"`S��)� �X�ݶRoޑJ��$�~2wi_jo�d�����I�K���5��Ң�^D&M�|���QfcK�!g·[K��_/�8p�<|3��q�sD2�.�H������f9J��5+ϩ�)m	��m�����&�v6�
s5��V/�0S�p ��)K׸�Hr�2�lK�L��rs��L�Gn��܄�d	�|l�$�#��6t�~lr|�w(�J�cvz��i��%��tk!�8YS6,��2�Rro��+�cFK�A(���ہ�=��b��u��1jo����*�n1 �1�wy�A�>��̽_��f�KT��l������I��3�u��.ڃ���'Im9�@��s?]�W�翹 \�z�p�mo���N��9��'��R��/�J��
�F\����5�v�f��ː>ɧ4�$D�-�������ze�@N���i�����-̽Ey׵1K��՛�}̷��At,���`�
"rڕ�]cs������G�,��,��k��1��@�}Y���lj�����{Yc�y@I�=�J�̱�'�~�g	i��7�Әt�S�}YL[T�Gg��h %�x�d�aO�Ž�]�s��{��=s燺�hGj���%����z~u�!t�O�D��+ّE0��~�����S����Q��s�I̥k�-�5�ӒhMfG<] X�$��W�����z�G���T���Pm3W��݉�i=q,�s����R��Gg�Zj�2S)2���4S8�J�b���:�C�|/�>��� �l��/��F�x�'*�I�PX~�"�^��J����HJʍe��F瘂���ρg�+�ģ�/0n�}�ֽQIu�l�	�3x�>���I�+^����U)~=w���0<���@X>��Ӥ��؞���$����6�j�{��Dt����YԒP��Y3*x>|B�{}��d�wȥ��L�iX\�6���͝�m���^�|%}���^yP��$m��V�&����j�'����t��ͯ�[+����l!�=�&���Uܼ��
Ĕ�PV��a�m��aMni��D�#pr��)X�fQ ��X�\��I�0G�Fym��+0�,$�I'�ӂ�l�8{�RP�{���g��a~	sH"F:8�]��;�x�2E�|{�B�m�D!8~ �w���-V�h�lt��]�h��N���8�ݏ�D��T����C�Lf���)Z
ƣ�a��K9s�$Ϣ�+O���(&H�DWa��Ś�@���m�2?�f�z�P�Y���vk#yގ2pl�g6I����Km�`�?�<{/R>�P� ��G��kF�ٝ�@���o�-�+m�o[�>��������RIn����5�)�R��HEs�/N�7�;�<A��`��9���O �)"r�=���XJ"g �b� ��Ц�i���<a�uxs�U��Or/�d v"f�yN0��T���᧚���Ք�5�s�i�S�`�p8����+�:A�Z.�S�^Aj\Rvo5�*f�����d[z�Mʿ|4%h��k�`�Fh�$Q�N��כ���͵g�`�33�����7f���S�)��O5RZ>)<%��|�@8bFOZ\��k{ڒ�����4<z����Z}���J�`��xw���"��8�y5�=��o9�>ĺW�{]�d�\��V�>����ƴ�z9�b�v�D��n��<r��nSn}+xG멎�������'���ꋺ��Ҟ3����x0E��]��n��[�r���	���im!�;_" �FJ�3�]��}P��l�WÈ������:�0����o�6���e�O|���t ��w��V�T�N�.�N�Y��h�r٥�Mb�A|v?��|׮��	��/�Lm���i��-�8��>�����ޗ�U��,���HK�)��tΪqe���$��v?��̳�E�u]�ٔ廜(:���(��:�nHtgs,\�0��'���
WLM����ф4�n�_PU&�P.) �#��,�v�8���8���yek�k���x5Ԓd��-2c޺�����'^zC8V��i/ݻ�4|�z�|�&����vx[�M�ԫ1^���o΁��g��&&�Fh��>�� �i�#s���`����FA�Ž����T̀�}6�j��]j���/���6���Ҹݭ��]~���U6`83��ٞ��g�Z��mDE�k9�g�k��yR�bJ�.���󓌥{���"賿A2��QSC�;�U!�Cl���7zp�|����,���VӅ3F���*KKmX��U��&�R�!K��*�S뭍��s"nsC�^�I����F�Ԉ��+E��^�C�%��������N���̠�QMkEo �A�`�v���ԩ�}�ԝ�S��
����v��;�`�c]sz4�Ђ���lB�V�t -����܂�X�S�m�?�˂�qƜ�ٖrl#��ti���)������eH�ؖ�R�x[p��mhh��Rs��K6W���W��y�Ɯ�+|g���D���q�w�xnͤE�}mx�SC��V�O��inhcc�p2���D;��`ˊAq���%���f���cS ��F| ��� ͱ1�!�C�Ύ�1�/;��(����}u#dK�
��y�-1�[��\�+@���`�ľ�xt6`ǵ�$��ns�b��������5��y4��T��/>�4��傀�۲�'�]D���\�?B̻�/_��jm�1�>�}(���S�$�7x�g����]@�>}����^��hq�v��or%7�R�
!qYy����x �[����N~o�?�^����ٛ�Y-0e�POߞ�>�"�W{,�g��.�ug��ѢG���{��l:A	��7l!8�b��J�Y���{��D!rJs�q$��	) fpx��xy���D�q�nܖ�6:5yT��}Ei��RB����o�v�	�b���]8O%�.m[N�=ܠ���U4.Ma��g̰�̿�ݧ��F����g�4�ضm/���4�h���"O�_��D���u�HDM�ȭ�����]�J�TV��%b&|{9�K4o�(��`�� ��h��&#�~�ٴ]�;sqE�%L���:?�<�ҺU�.v�u�ǃ�#FjbJUp�\�K��U���ؓJ�h�
Ե���v��y���UY@�xVj2]��st��9��02���ϳ�4�D �cy$�
ECBn ��@�����������8̾���4�o�Ҹ���4[X�M�y��v�g з����}I�3��z���Q��/��9�'� �jɕ�[�ԛo��g��5�ǆ0��,��
��B��ÉQ������mPe�D/CصJ,�w�Λ\����o��bV��v`!�ora�U|�DV�����B�0�g5݀�)�`Y�$⥩F6��g�R�3ZvyO�@�Φ)��t�p�Nˬ�7��WS;�{�T��˰}�1�5Pk�b@����ݠ
��ì��|� م+��92*��b+O_VZx��]�153G�#8qv|�l�� �,�2aN����# �.�y��E�W�I��#�sx��D�5�vaݺ�H����Q��H,��>�O�ؚ���OX.���혾k�w�L�3@����0	��p||*�;��y$Y�E�!].�\���,fx�bKEK��"2?xn#(��-����ʍ�ã�3Rw�Й�#}��������iH���L�غ����W�ߚ�s�&��M��ֶQE���V���dA6��9���~�ʿ<e�EQZ�+ͭF�g�'���Q���u���k3P�Fŷ��xY���Z= �%7�G���˴W/x!�8��lu='�c�Z�h�m@w�����8ڝ����\g�����~-����}�ؼ���%ڕt`����'�~d���Q"� W���"R��vԠw����.��䈈i�u�`�%I��l��1�)�X�<U秅u�@�"�:�X��U&�fg0����VG;QGx��w�k4���3�9�!)�h�1�6��Y&4��?�ƍy�u�(�){?�wx=�����v?}�a��槈�}��㎜���-����r`����h������p�S�m��_L��1��&�D�:�R���{�]�D�����r;�E���'�HUԼU7�@���sh��X�8��\.���DN�Dt�P4�לA�&��L�'R��&_����%��<,,
Z\�b��\��._�[��j���B�\&e�=�L��&��)���E����QFh��X{׭��Pn���s��������Q�o��7N�%C�C�B�dy�<C/�=���s��[PE���[u��b^V���Q:�-��ok���ʹ<ю�zMȑw��[����"9������O���Q��V��9š��{91(w���1��>�����k��d)~w���D��0[���N�m����J�K/f�;�7�����H�rD�ɺQ�O�\��(��R}?�zb�*<OL�f�=�P����]�e�ڕ������Qv���0^��@y����f��5G�p<h�v�Y}�.�'��V����r���GAS��l�(�ODz����5��mSsq������w�֥nyC���Ns|a���K�?E�ϰѩ����-f�7!/�DH��9E&?�<v��l���0sB�x��~�6$�]�vs��f��esyXн�b���VbP���?ފ�����������?媢s�{&� �^z��V����裋i�%��a��*Y�E?�̖������+Ȍ��O���4fj����+F��^�Ts��X����C�T��C��aT`7��(��;��`.�S~�Z�poE���tݷunD��ӱ"w���ǂ�ȓ����Ei�bZ[���!�Z�/�цC�D�l�h��|�{��tS�IPH����?������ 	���8,2�#a��L������4ͭ)lX�t����R�|f��&A�W����k�����˃�1�[����"t����ߗ�����ޟ�W%d��YJ���ER��Ι9t�e3H����/r�eUjƁm1��$��N*�Y��p�.:�
c�7ťpLߧ��jQ���ZeV�,"t��ٮ��=e�/�-_)��n&_=��r ���TVJ��m�����*6�$p��5fw����] 5UT�ҙE4{1��w��F$����Ǘ�'_��:�
<VH���'k�eQp �qx!g����*�/ �!�6�6&H��_�3�[�P�3��K@Q����"Y�]p�L�e���u�\F��Q���-�[�e��{�cȔ���Y�|�E y�f��O3t!��A����ūB�u�C&�[���J+_*���H<\~~� ��@^d�ɿ5��G���xoL�TR	 s�=�LBf6�dq�$�9dE,)��n��N��r:�E��������٢�v�@x%��[�����~�����Q\���VE����ξG'Tl�+��4�|���9�(HpT������(���P~ M���-䜋��n��ݜ��SS�/���3�����ǠϨ����H����G��|p��¤/0�P$1I�=ɐ�:_���]�-;;�ܷ+i��%*��)�K�Gs��Ny7���=~��.īy�'�K�d3:�wr@��_��e]�g��Dm�mh�Ӕ��pK�����7��ׂA[�b������D���(?d�x��n$���H��$.��0��Z���2�Fh�߂'��Ʀ��U�r����qĞ_�'X�i�~e1>d����Ka���,;O[�>�e���?_�+i E��n�K�ZV˸�����=�����t���p�i��rRʹR?$*�%���@;�l� ��7��6��x��my�ul��G�=&�;]aSz�<^��d��	x�b"���obϐ���!<����Y���2}�����/�~�|����5/L7BHtD~X��h^}����/3Ib_�z���~���&�����Dw�:�Q;��9s"��xF�ӵn$���v�\l��zB�}%h�Ф����!�0eӔ�luMY�T�a�裉�\�p ���]S��h�.��K��"��ɖ�&��џ�*:!��n)s��?-�Ѿzb��E��4'姈�m�ϴw���u�[m�5�0��>I�^�=z�S'\ f��/�V�_��!qn�B�d̂�,G��>�U�ݳ��wWd�p�&cf�����݇ta�Ȋi|�����Zy�q~�t/�M��4֏��D�ܡlgP3#S�@Ƃ/����;�2� ���/=1u힅���Q�(��ά�:JV����G�
����KIc43��G�����,���6��Dpo!J��9����T[}h3K��-����j&a�T�";s���LS�7 6���ֵ��_x�o��~��P�d�R�׊�y�'9G�L�ᛟ�r��j�:�8�=�" ����fH��Q2V�@��������6`�/p�'�nQ�i�ʡǹ��n��M"x��{SXcܓ��3<�'؃ẗ5N�-AA��ujB�2���u�(��h�O?������D�"�F� S,��� Tkv�P���+�li�3�p��[�ǻ����!��31M}��[���pt�9Ϛ�j%o�t�o�{�p@#/&�ݝ�>¹=!V�b FL(ݜ���݅�ﾷzwgZ�9�kW ��A8ڤskbd��$���ɟ�A��Np����a��ψo���2���K��	�����L��� �d׋m����:����Q�Y����S	�3@�{E�$83s|��� T�>	��n���:I!׉��Y�5�#�j� �.Rv#dOq7~a{�v�Y�C<F@�;s#4>u	z�n�	����8�=�Ux�_%�237��wϿj_ؔ/���[�����P�i`�e�9KdObϼq�n�� ���S���6~n�`���W�T�N�˸7���s�?��0w��fO�7���Xֿ��v>Xq��
_>kZ��v�oأ��b���i�cTvVZ�͘m��_�KUߛc�=�N�$\Z4�<�����C�z��Ue�3Ce��S;x�fOZ������)�WU��޿9�<0�y4���hK��^&�O��8��`��2b3#�҉ƜG_o&���d�@�M(���*����)n������aJ�{j�_j(���i�H�LI��?R�k��S���u����U�~���y�Ŭw�ᖓ�b>X �'�V�1�I��{�������X�|#H{�5�ʧ�d��z���+�m���복ƦJI�����xmRJ� ��z�����/N�5�jf褷�r���� ��NvT��
p�O.��Vz	����#;z���H��;'��6��wg���Y��SlS��>Z��%7<��xJm�x,��@���ZD�Rbw�p�Ͱ�S�SR_=�ZH�s;x:HD���`Pϑkq�)lQ�W�"/-��dMJ|��eH��1��[sO�ӟ�(=zy�A����D�:=/�v�o�pP[,�Ք�9*ϭ���<��!��V2�[�����kH"��_�Yy��]�-��1�/����ϖi��f��/�M���4Z~Q^W��k�Tn�۞Oʥ���U׾�ش����Y�!��i�2W7�����̮j�5/=AwAL[�W��\y���y���J�MoKD}�9�+�����}�A����r>[	I���ln���ZYL�m9��ӐW�/}�0�w����Y���mt%�} 0!1��܍���u�x�$[�Rx-Cj�t�%a�zѹz�_�e@z 	�P���][��q�w���j�3���Xn[���t������+ tV�+�,{�bQ���Ǥ�����ζ3���³G�!�`�~z4+��}Qꮟ/N�Lq �eֆ'�!{~3�lO%��X�h����DP�����F���Mk���z��c*�Q��߉&�Ӛω�ǧ�4ɴ\8�`֙��cӐ�0�C��#	�n�|����7W6O��z�O���O}����j��Y���F�k��끏:O<:T�{��ػ����
��� �����owl��wl�/�Ծ��ߊ.�0��<Ϥ�{$X�*�2��+_M�bk���ύ
bIM�KP������Ϳ��,q=��>�e�!6��7[�c`�8���f)
u��f��Np��M1e�9t�8�L�}(��]�T�$F+#o� h%��Ȑ�yI>nF*L�^ͤ�[?�7G��N�.>�d_�<D�`s��R	q1��vm�(1&}r�実��~%RkK(�	�b���j�2ѭ�
�H��)�FQ�>ZA�,C4#Qb�No�nU��p1�ҿ��̮���7��&�G<=��5�[V����[8�����:���Z���t��!��Kd�s��j_�V|Ʊ7�J�[س��`��Q�쀠�<0�Y�i��-�/mʹ���5�����^��0dǝX�����	�7v���*���ob,D_����/E�u���z/!)�ܑ��Pi��p]'���⏂$�t��v�b�5/��z7b�Snfoh�uO�s^��)��;�ؔ��o����C��S}%���O��J�iW���p+��̳��	�佚v"+�W!�$[���e]kF��z�[���~�f!��.ň��~��Gި���A���6�b������+�X^������B�;���M|L���8r������8 *�o�3�q����^�'�2�W�B׺��"y[�aZ��D����s�D�� �Tu4����L:sP���!���^%a��x��b��ǆ7t���'�IV��.4����P��'\^��Un�����10º}��N7�9=�5�:q.��8���.�j���W-ca�R��;+ɢ����.;LR�`�z;/3B���";����!�l�et��g�Q���cp�r�2��F_E��Ww�A�Y�_\�lG~h�����#8(L
���|�NBB�㻗E��zۛ�6/��~��pW�Wm�2"��Y��).#�z�?�8ToMn���'���I�  ^��ƆG�c����b�o��e{�����x6�N���k��R��u��
����CޫM��2$�t����d�ݹC�l5����rR�es�eL8�;���j���Zr9
ڭ@������Ǉ�:���wӎ���1�e��I��#������.ǽ�7�
,}7�P4z���l=��܎%�-'�i�^<�
K ~>=0�� +�J��Fq�b�It���|�0�V^:�2���1�/���6��j �z��ή�a\�2Q���~e#oXs*&�4�S{��4���CG.e�H��?���ߚ��	)�K'|��3�쿼���)�������g�[EUCe�����4'��?ǲ�w�z��:�H�G��c��E����`t�go�yD�1E���jJ��m�$��'�>{m�(D��bY�%�bT�c�
3�81�/XT��F�j�oL}UT�&�I�$��Iڹ �C^s%_�Tj�mp�8���'Z�4q9�"nj�.��G����b�Q"�s �v��1�-��������|kB�|q�	m\�\D�#���
Q���T���N��ax��T�����*bo䋇��z��3�	������`t�ɲnh�o�ʡ6�ۊVЀ�[!~c�d#�� ��f<a޺���|Tj���n�������}l?��E�������h؏�fJ	Z`���]�l�m��m���ͣ]�5<5R`<IWW�*D��0(3��; ��uv�\�ohb�0��L����3
����]/	;��߭X���h�n϶j�H6y???������n�O� � o9J�?�c��i�M,�����r���Q�N���������.>�
��#�|*�P.=?�)���[e���Y�o�?�}E�#��?�_�}��"��"��!g�c��|��,^��&���r��w�g�"�����G�b�A&G���w}
�G*d6����h� \g!q棽���H 9���J��v� \1�����<k�nC�>��K<���t����u�x�@1Jr���Ƿ���gN'��W��J�},F�y=�Q��v�;22�HX�S�����=Jj��%#������G���P?�ɂ �3����.V9�����T���uE���F�/���sα��T�*L��#���z������/�U� ��B���m=r�0Uڋ��_�O���ى<��PQV����ڪY��Q�T���/��e�~��]kQ�_�B�D2�\�B<5�oiW �-UKW��-�~��=XX� ��T>.�bQ�����r�+��]Ȭ���-���_�� .��5Pr=����$���-�V�A�o)EڌQ	Ĭ1kdR����~�&�q5ҏ���Z]]FɌV�oE��7/�_�"�O�<6]T����
؉o��g ؖ��3<R?�Wd�p�mI�ߝ~��]����\��=6DZ��鈾���%Xo#��)���J��l�2n�̗ܵ���u)�c�SVE˶=�����ہu:z��f�.b�����-Ў��?����΁�ힷxU����)6�&�)qm�s�͝�h�di'�7(�y�݈�;��N�N,�(mp�È�]�j��)OGgt ����=6(-� �����*o���S~jIi���'�w�<�m�i2pj��s�P2+ИVu�uh����>Aڦ�y8o�� �� L�qw�޺�_ ���`�r#����NT�.���Yu����������!.z6'a��K���O%5Q�%a���Tr� .���QrRM�P³��Q��ցg>�ʾ�b�"�D��X�%�d.�l�RO!��۞ir�W8���=V�/��(7��i���6x1P�Ѣ>d͟�]$���v$�Y�fy;C��@�ٳ���Ka�>}?������
'�hS��D#�wn�'�~$U�����e-��w���m|��ev�`���@ڷ�ͪgH-bH-��+�a��bg�q]�����ى}$RtQ�}��C�T�=����J����h��z63��'���s�¢R��J���)�$}i�,��;|��Y8���22V-�^5։��mAds�=�/uG'�*�)%���4�]b��& ��E�<�}*T#�LaaTN��_t��k�ݰ�/��u5�(�������N����,��0%�P�ښ�$rLt�af�R)~��r�{E�y��]�����(ѧ'kҶ�":���a���sy�F�OwG�w|�)�@�T��Oho�x����Fݢ�-����5��y�<�>|ͯR�}����*�L��l��`~����v�b4��p��&���1斃j�2x���c�R\^�J�-�T$'���f�b��w?�/��Y���p�Y�2n]2yދ�֮��'Ym����ӫX�&8ŵn��A�������:G�ز�j����$�B�m�ˎ����+벢t~>�XP�<�� McM�'�F�ʽ0�hQ�uci"1N���qrZ�'N�z'�$��=nI�f*���8���	�!!`NE�*G�/���͕��f����0׵̛/�!��L�qN����#�,Y�/C>|*5P��-(�X2�r,���%��lՑC���ٿ1mr 
Vj��ӧ�H_�fmF#�P�k\�u!��|5K;-��ܼQ7j/��4a+x��t��X~��3kI�TӳT2��Q9(-����t�Ls���1CbEX;e��Г1ҧ�<�e���K�����P[��\���b��Fk�e Eol\��XXY�2By��$K��,sʶS�Ĥ\��ݱ���Y��Y�������bA��?��:��$��a�ּ�!�DbcV���~����Zf�\_�TW�\����S�W�na�]ʓ�b��-�D~6[��9�.�����n~�@��G>!-q�����V�|oW;���	��a_P��bc�Y�d[F��У�b�8�� F�՜�q>���9N=�ke�}ĸj}�P��g]�l�ݼ956�A6������V�tUN��&��|�$9`�(�;��V��PY݇Y��� 5�w�}s�RQ���	f/ ��1f-7y.���V~ʾʟ�\�n�{�u�U:��lD� 1ޓ�� �l	���[��38E]�O089�jԵ^��]��oIsx@��w�}����X��ŷɂ�Q����,uN"��/��鹟�ۈ��# �mF�.to�T��|�zo�G�%B㳜F�~�s}F�8(P�����p-�����&����n�[�к�[�B�8T�_�z�>��;��ƿ~��Uu�W�(��PAx�L,�����z�C���q��:L�E��9>J�n}���$.������ej����՗��po6a_¿k���kj�/�WPGr�S��:5;���������f�%�#�E&g(h��}-8[��Ă{e����kb��C���ݝ�rmd?�I�	�B��p��zf>C��5Ie��*�V0=��p������t���
W;?��D-��2'/�)�Ȧ����L���Q�1�&-⾜�ԇ��q�(B����1s��+�j��i�Z���y;S��m���
o�N��A�S8��_�WcI6�B�zj~������f�ɮ/�ZzLɩ�LQ�(��l�R\���|j�,��;իK�
��@K��:(7�Z*��C:8��4�̣tY�]���uFN�p0�d]J��#?_*W�;�f���m�nRkx߬��x�Q�d���@����ɤ�7I��ݑq��};F.�
���[&l�閧����>#�`�n�#5�$���K|""4÷�wx&888�777���-����
����>����ă��'���k����Z����9Wk ��-i��6��c��K4���ܖ�K���d��Xb7|����l=Lqf*l�s�
ط�ܼ�NweY�/#�c���^�wv�:����HrhJ��Y���(���~�s�-�(Ҡg��x�.�HO�5?SlJG�@Ŷ���,K��S�~B~�e�`ϵ�oG��L�H9	>^��o'e��B7e|hz��o��(��b��N���D�@��v=)N�;n�lծ�L���81J���O�hb-)GuD~��nO�����V��o'b���E��3�V��)n��KKw�O�{��i���\��(����ULp t����<�J_�,z���~�5���yOZ�OG��ѯ�
\E���Uht��V����
摃�]�ł�W�ԫ�I�)'��C�mx��p{������y�[�*w1�Q�dQL�4�i9�+e]5·�Sz	�"2�,��/x�8�Ŝ��$nT��
�A;]n�H^��ЭQq�`�	������f��-#ae�T�d�32*�f?��>-�C��x�����dR+�����e�t��)�;'�2��NuY���;a襚���#���a�9��'̛m}:�X�Uy�y�W{�Z�ŧ��
^C�I�e�2�:�� �=�K%,���5E��H�K��3H0�'-�+��!XY�iV��?�u*b]��p1M���(�S���1����s�79͉`��/1��%J�r�Sh��kGJ��<1��hcG[]���k2�+��0������ʇ���˺O8���'}	U)>�l79H���xU���+XG`=1��ל?��w���u!���G�Y��c�./o�(�;j��{E|[7��+$6�a�� ��eK׺�"��M�"��EeFb��*�'mL*l��/�K��C�[7�;A*7�cTD���� EE�3��O�?��=|�o��-���q�Qt|��j��-d�%'�1�"�5�4��gJ_����O�p�y�<L����z1ܦs1�����f�^�σ�)��+,T�:j�*jq���҃IwK�ɭ5�@G�v�4.�H5��O:G��T&���g>Qg���Z�\'b:����@@��fD��6&��zk���bY�O�	�	����A0U��K�YL�}n���\=-�����%�w0�bG��&?)������j�U=UT2�lS$�Z"�(� �xR�.O��R|��60K>�⦰�+2����~e.!�qpG��.�S]H>k�i#��䞽��fx\�zn���X�a)>l
_�P}Z�W�Rǃ9�W���RRߍ��'y�GiV��ʚ/����3#��}	�n��7c�ZY����u#�S��?�{u���v���ח_��6ے���Df}��-�F�J������[��%�#B�GDNl��
�uYfMe*���Z�U���L�p~Km- ��٥�"r�</��b�tgQ)>fL��mE��@���Du��u��5\U�u��y;b�oCc�F_����{��m���K��7�Q/ �'`��t�W�����:X>�-���_�V�f�������O�RN��"�5�"�����˒�ڧ߳�e��K���~�l5�z!X�Ć��ВRBl@�Y��M���תP|O���������Yօ�����Cpw��Y�!www'	����m}��o߳�s2������Y]�T�SsVw�j4�{��LJ�0�G[
�)�Zi��g1�N�i�#���:�x����!����W�a씬���z�y�]Jc�]!���~�$�3��/d��z?h~����q��?�L4���^�c�<�c�Vt�X�д�7�w至�S
׳��O�Y;ԩZr��sv׹9�h�kN��h�"=�z3f�vܠ�7�V��L�{R1���3�T�t�f�8��â��|�~��%�1��fg\���c�l��6����<9,�,�oG�&�l�u��ڷU����������ƽlB��݉��_{���K�Cm��$cj��M�0�qwF����oL4�"��;]�����%'����>��`�6��	VNb���Ā���MpK�Q���4^l1��V$DW$$�����'�"$J��_��Y��]�[��|M'Im���1�<�.?�D�/��HvZ"<g�� :�fE����-r�:��ϲe2%ȏ��m��t��q4�>��w���,�mL`��P�����5T���$��|��zb����!�6�e"��~�JU�р����i:uD��^��C|���xX�^M鬇��t�|{�4�)z�^����ZX�s@����>pt5���%J���SLh����7����܈�K��2�}{�^;��F���V)w����¥y�T����t���)su�	�D����B�V�P|���v��'��x�p �B[�V��}�RN(y+n�'�;U�g� �F��J"$K��ܰ��$�C�sJH�e����%���T}٠���I�3�o�h�����/�~��P�H������A5XY��tOƇݍ�a%���@��q���qN���Wi4��2����:QW�0
�c�u2��s��z~����B|�@�K����C�2[� ����خ�� ����s�%���P$h/�ޤ<.}S�|[ �^����/Q��N.� ��ړ�	|L{R#��S��݃�Z�I3��]�t&[ڜ�[���:��h딀0�}����l�}T�a%��R��JD�M��c�i!T���1�|�Ce��M���:�p��� I��{Eİ<��$�؅�$���A���(�P6�duR��?P8H{p�zb6e���vF�V��������/���^L|Py+�)����>	B��͈U< � ����9~�A�������G�>�;Iߵa_��.5"H�=BI.���Qb��EOD�N 0�#M���K�U��"D�O}�&1���\��a��k���$9ˬ-��<AHʤ/��
C�nH���5+���������!����5��^���mW]і��t�z�m%$�Uނuٲ�����":xŹy�33 ��/�5.]�:\�v�,ȳ`��z���a�ZNH�씒Z*�n|�n��:��,R�<G�?Kc=���L��w@ƪ�^ؐf�:��b���{���*v�$�>��	����+t��om�m]�KpLZ��n����t��<�Ä�ӣ��$j�s���'~[ˇnc� ��B�{^�.�u	��뜮n^y#��͝|��f����_@�v�s����4z���� ���<&wu�^���H��a ��ި��E��`sKa��}���G��~�.&rz�l!m/�#���6������ I��.�<=8x����/��)����Rպ�+�v�k�:��ġ�x��[��]�o_V���ؾB��C+NHD�w�%Y�С�)�ن���O!�ߵh7�i��Qx�x�׎��;�T\���A�"Zb����*=HX<��gB�0@c���5��,C]�����E��kD��1Z^�d-�_�,�G�ѝg��1ڱ�X{��+]�j�P�e-yZ���[je�HB'��i���ᤐL��xИ�zv!�}��e��H�ǟ��|]n�G�=�^��&��*�,@h~Lso�<��.,1�=)*�v�� *�1-4wL�[�;�t�I�������� ��;l���%Y.
-l?��C�6�܃�vC��KH�C�^��8巰}���.���ӫ]�K9�q6R�D����%]g����6O{��_��,b~9���N�����C>�?\��>������-��%%>.q�����q$�e��]�����U|&&L��$�}����"��u���v��b�R���%U�����.��+)��2AE�j>���u�4�-o�|�_rr7?f�M���$���0u3�����p��]�4�=A��'�V��_V�K�J)��\���������d�ja,b<�P��FMɻ��`MS��n��=���N� m��k��pD���K����"���P��t��5V���n�(f·��<nit�<�~�b��ӯ6��mt;  �]�V!݌ۛ�f���N�[k�( "yo��_�;=UQR�9ل�3��z���{}�Q�l~Y[ԥ�C31���|�`�\;JG���"K�{ψ�C������9������3��O%���t�)Vi3�#@|��R(Wk��vJҎC�J�v�E��F��'�����iX������a�ij��Nl�-�k��N�� E{<��O����/\ļ3��T�˖lHқ�+�i2��!	�7���4�׍���"̡"�5ж�0�?1��Tf�ģ���Y���4�5S�H�,�Ξ/���hS�ab�E���	�J5F��Ag���w>Hu�
�?�-�ߘ�=�
ӱ���z��Q�e�%K���F�9��y{�@D�����md<Dy�g��l��ba��#���[�V���(�7Y�A�����k�S��Ľ�)�Б�k�S�ZƧ0/��θ�N#�Q����f�/�?L6D^.?���@�'���Z��a���N4����(݇����_�fu�:6/�Gim�<��(����J^����|����^�B\�����/rdj��/�:L3ܹz����?���U�t��GYyg����i���J��ٲm�����������!�E����M�Slғ7d������*�7G��a�t��{#���Z7�,��w��Zj�t�d��#�:(�ZV���i4!�JVܷ�y�W-(���f�+w�.�g�#R�As�9����뵐����<�?fi��hi�jtӬ�}�XX�|���������'iX�}�I�	�lX�+��;�Q�U5�A;����xC]�r���&\ޫ��Ö�ˆ���'Y�k�ۀ��d��!w�����H��u*c�����O��S�0��v�t�]��n���ZӲ�AT��X�]��,|��LT�b���눃���|�{Vy���5[�������!����+�kM!x�#ٕ�L�{/G���O�h4�0ݪr������j�<��]
�o����R8�n����tX�a���J&wi���f>����r\�S�Uo�l��R.�,�}�w�i|i��1�V3�x[�/ͯ�L{	�K�fR�y��1h�"&�Rb�oH�$�>�&o����� ��zf��'!]v�S#��)�A���3:�_����j���
�0�����\"�h3K���_:Rݭ������?����:��ٕ�5'�ҧ��}�:P<;ލB���b!�->�p�U�+�-!��c�.T���dS���|2�z��k�O�Du��!�!�rK��Ԡ�WM� *I^��Z�����S����9�-,I��<�e?i�$�Ϊ,+)��Ǐ�kӷGנ�-N�W� ��ܴ�{0j�z�Vn^�W���j(}V_�o���ʊPTꤽ=-���al@氯7�;�!������N����z������FP{�Ѿ]]+�wZH��D��,��_�i���b�!�e#p��}���q���X�ƨ��ud롢u�������QZ(,͹���O��F��4#��A2�f��������<����yvt����y	��u��$�s����es�'Ǜo�[U3m���V�/^��^t�
���!�$���l���P����5X/�jl��mm����y���r�0�{>б'`���O�R���:p���������M�w,KJ�~z��mۭЌ�u��ظ=��N���} �B��y��RU�uS����ڝ\v79@?ܓ�n��Z���f��o���h��O�A�g����W��֭FmF�������El)�3�yT�- �n(��#��Xr.-x�R��Z��4��>��<�CU��5���SY����y��8�"��L��"�o10�v��<������� n�Y>�L��sI��6��4�mCA7P���ZU8�،�Ȕ7�M��<3|8�h-��i������N��W��8yݯ�]�P�L��bPچ����~͟a���F���Q����@��D5�����uT�{�abXS-�'Ŏ-[6�ހ`�q�pR��޴V�����#�m@EgJ�M���"����.X��,~��2Z�2��"*tv�����Ǚm���c��O,C|o9s�C��S�F��G.*��9<L8���:<��k�ֈϵ�.рP�^�f�$��l�	o�	����bT�C�T�`�
����#�n�EB�Oll�{���xdێ	y��1?�R��7��uuǰ)[/�_�x�	}b砐�uJK����Feb2]pǦ��<~�O!W�Ϙ��XӺ �J�7r��h�b�O�,��B\j�"���M�K�p�B�+��ϢA)��TɊ8I{lv��� $��*�dȸ����ō��ߨ��<�ر��Y6h�&���-��\�*�
��UV��u���L�sH��Nq4>��A}=��4����<pupA���	�4�;z��ڈq���Q^�]��,�N@I\��g��0⺫p�H�ڟ5��<`("�f]qØ1,1��e���,��1z�H��'�t݌%Q�ԈI������S��e[Zȣ�|9�,��H�-�����7[�QT��j�P0��,ZZ�2"�q�����#�^�G�u�%5��3y�f�i
����i�t�߸lތ/��4��f�%DJE��hJ^wy]���Ѳ��#	fn�Z���$��Um�Ł{'�ج��׹���2��#��9Xk���V���p8ȿ�AV�Ծ�a�	�#�h(ߝ^����K��y�9�$����Q�X^�pV�ٟL�he4�v(&D7� �(����+,�e�a Å#ƮB�c�N�A��ɯN��T��Mv��RP�.�9��v~�sJE�����+mB�
���3x�G��Ӑ�M��ՍB��I9�)�f/X臬�jU̞�f)Ǹ	>z��/
�E�,�k����ѤԢ����uM�g��:�4J��O�&��m>�s���m�ҿB>�'�ja~WDy��WP��%�|;��5֔���R);�[k��>F &ƣ'@����?���DRg_�i~b��a�u�fl�8��kp'�c���6�{���HF��^u����C>�	���1h8�9�|�����q>��yvS����i ����l�>���[�$�
��rll�G��
95��MTDb�����XYQ�R&e�2��bL���F9T�+�r���'{�=�FI/fF}�b
��I߬:FRe���T����\�rD/~������^��#@�'�.C_�LAh�B!�c�حk��g��[/J�}���B��*�7��jRmz���.����f&"�46�7
����EE��Cm��*�U�X����<�Σ�8u��1��Jgw��7�'㷁��;ӿ�_Q�W	:��f�2g�.J�\�����׎�:o�#�/Ԟ���.So�0����C�}fj*x~~����޴0�wy"��wt�m�G��Bd����T���7Gji}�W>��q�y�:�4ݢ� ײ�w�|�������0^&�	ʅ��>�ʥ�U�B�#b����@L��U��C0�h,��Ư���/E[¿S)nw�fz�[��[�v�g<H�s���bi�΋�Ƞ���3��q�F��v�֖�"M��	I�Ю���bݞd
xK�����+��E]v/��v`_I��H}�z�f��>@��6m�����#ڰ����*fJ�4�	�DB@�4���T&b�p%�~�����%VDp��'���ɯ�d��V�Γ`yAue�������-�3#��F�	7�p�����D�y��WG��ja��|�Ҕ�y�����w9��Ӯ5����r�t���b�*�X�L]j$#3XQ�bU�o���xC1fO��?NР��@��v>4;kR��\�ˮIw�4��f��l�����ǀHÆȈ����k��y���
��u����Uw���X�<[��;"��}Q�bO�p�PW�'��m����^76�3tpB
��o�n;ÔZ#v�#Mn���
����>sD��HqT��G��m������eD��Y�Oo*�͊/R�uW�h<����t�/�������l�!Қ�ua|�i'�ɑ��q�)l��Rk�����=ٍ�4�8:B���9BU��g/Q�(.�|x\�b�}�Q&NJl�S����g��&������XC���8;����s�.��}�"H�sJ|�s�g9.����A�%+��I�Ŏ<X�|@���'b;���������/�ykAE�*�&!}jf*��l��
#&�����S�7d����"��:�K��?�5�2ѐv�� ��޿�s��(
�x��Z����p'��n�"v)��)	9t�9��W�hD*��%�X�w���YB� S݄�K��N8�&�,���T��?��ߙµB��i|�=-z��G�ST-�P�b��K^��.~��.t����ݽR�����Q��Y<lʠ]7 ��4����(�{��淐�����`-l4��=�*1]0|SNIm�ޔx��Z�%��Ig�_9���|�(�N���a�|	g"�lF�󁝸��u�mEBk��6 �86�a�Ca��ɩ�3[�BEaB+���� M��п�H���a��H>ЕS�;��jp���?+�֥w��,�-f�b@W��!�:��� ��%@s��	X�?i���5�E�Sa�+9��-�S���-ҟ>���X�뽁݁�lQ[�bɭ�!��罛�o�������д��	�>>�Sf~҄D���ⴓCc(�n2����kT���_�("zֳ�����V4/o���yٻ�������7=��	���Ss���i��E�X��#��i,�!bt�(����SZ9�m~c����'�Y���q�j�QZ�H���q�sC��М�4ϑ�ww)�����2��ڠk:v*�sM�������p#B��Jl��L�����mZTL{��(B�`ۭ�" [��L<h,�>Fj�1��xw\�{V߰���o��G�B
���w�-y�Q�I��2��*��LA ��쨨�$�C���}�m��zX�|p<��v��A�zh�E?�������ݳ�I~���p�iM⨨�fGA5p̭kR:X�Q���,p7r[��#�Q-�L�bc`�Qj0�<�h;�G<�T���(���aa2���)�
z{}�ti{�t��x�h�������5m��z2�t��1R�"r� ���I?\�я�s�P�� ^��.u8��x�u�l�
���t�:���7��%iwQ�B@�bC(�:?s
�� #L��  �&��T"�k��Y"�D�vzs��&q�M.�=��b<f�����P$\�����>0[sZ�fȬĆ��_�kG�ɇ�_�a���'�<�O{�m����7����E��G���=�̰,�@߲d�T�p�fg����s�<c��M�l]��L<:�}k\���������֏���~�'	sz�{�K���҃�W���v$b��7��߁h	�<�!$�H}*�H���,�%{�<c��tO[�t	���5�����Ǚ��_�I�~	��ތ.F�Ӄ����$ٜN��@pM}���	���c���ݟ�޾V']U���JٯKOT����0��!&S@�MIM�iwظI��?f%�F��l��!�s�l�.oϣ�㿴�3}c��()��VռMB-I���s��<,�}���Z�H<ϣ�4u-<;>�@U�����u�^�yą&Ox��븞����z	u����C�1D���$N Ø+����n^�RLbշ,b�p���z+ ��̡>a�f\��s��yF�����?�?�-dI.��	�T�F�VV=��q��"�Y�R�v�m�R�RͿ����3���P�N@����u&��t���X���~y�[c��Q�cp!c t�4z��Q=���-��2��5vsJ��	s}��N뺰�5�hq�J�|�1�"�a6�8l���_��������ι�j�P[��x��g.hl�"6�������c��O�@�KVx1s������;�z�@�1��@��W�	�܏�#6���ZRkf+칸
�r=����2��\}~��L׷��&��(V�I�Z[[g&��������1PJu'a��P�0��k��y�p��L|���	\���!/����(����������O�Πu���,ϙ|d�9��RM�c����ȁ2!j݉ȇ�_յ͕��B_e������]��ҥ�K��kl`e���G3�E�B�"J�<e^O�(e�0�| ���1�N�[mqU�@�`$6p8R`�����6��M���b˳¬��/�{C����J�w~�k�g"q<e��I���F���9�.&� K�w��M�1b`�Xo�Pw�J�~lUԧLE�|�ap��S�H��IC�d>�Xw�����H��E�@�����<%c;o���(����3+k0�^�2좻�f�s��?�.�KS��&�W�o���W&�$\|�GbjQh����ԀY��d��+TDkmQ��q�^�\��G�U�3��D��_@d�n��e���������X3&��Q��D��x��[��f��� �Q� ��Z�� d��C�i[���������QN��l�����7t�	m4�Ӻ3��Y�gg�ry�J�!�S8l]2�+�0�p �L�z�����I�Js7�"I��]yg�NIP�;$L�M�VX�����]�n�^�ueJ҃v����zg�K��{���SɘcE�`��vw�8�o���<R�=1�^���f�=}�m.77W�GlffvF�h>]�&66������"a��[Ss�xq��,��ϐ|fV���Z��Z����|~�.#��z>�v�O����c,[�1&���Uo�D�;��Nr��vV�3���.��W,{.�n��&S��2��3��$��:��6z�c����jE�#c���@��~����L ~�!810r ��3�]XT�DV��v76*!��W#�VPW�s�z1���|��Z9����d�$w{`4�e��_c�p�]�m�Q��fu"燨�����Y�@ +�H�a�8�O��!���!*�ӳ�G�	�k�P�\asm���.ؖ�or����8��1`IN��7�8�r�T7��з�3j�� ����"�	�����u4���f#����bs�����y�u Ona)C�ϔX���F�0箹B�g
�li>��& ��f�us�t����/}*X0[�"@NI#d*�?�n�1����k�o��Å�nN��(@	�����w" 4`��x�i{��݂�.f� �7��n���D!���_2�̔n�)'��v�/ՄZ"�<��z{����˩�8�i9�L��A*��?湊C^Ԩ�\ߗ�_j�6����j_�D�vu����C�ˤ���Q��l_^^6_4
읜�҆���d��:�>���5��p�dtjmK`n�n+�P6٩n.�hbW�,����O���ƵS�d�tl��ܪ�Z.��SR�b�WIw|�,�b	�K�������;�0]��O���]���5��<�I敨���H�ϐ 7&R�-P�Ҏ��?󯔤4�)23��9w'] �7uVi��uu�U^�- PNM��2�7�Z1�j�ڭ�Q�w��Fx�#(Ä �� �[�>���|3f`{J)�@_���\�Va�t}���J�RQ���*�!K�s�x��e����x�� JO�}KIEB��s��ü�{e�3"��#��H�m���ۉ�H���~r0�- �g,Ӎ𴒦?���/���G�?�Q��*�ww���ca�@,��6i��yh�Tnߐ	
�S_CJ�=3uw�|S
��zm�#� ���SVd4L�hvV ��Z�ʪ�vo��CmP��}c���Î����y̧Nse�� �&��� �߳��^��_;�9�O�q���z���d�S{��Tֹ��WCעi�C+F�$�x�w=&�Iɬ5�O��j��Sq�]�ӽN���0��oF���-~�.)�R�=%rɄ�R�#������3�$���y����P�^H����ʱȑ�D�,,,�_>�}�V��b�E}�H���z����t��n�Y�5�x8U�_ƶ<�#��.��
X�-%'�>8���p�M�X/˷����r��mH��B��]���3������B�P����z��{��,��*�|��w:���Y��2��S)F������jR�	��f�]5Q���@ ��������'M=�6/; TO}��&��\oY�v�)����g�H>z(ǯ�d.GU�U࡛�f+Q̅�P��(�&���S:F��vMڦ�m:� �ٔ�jޱ�P��*�lK��z�f�n����_�㨨0b� �>�����-���5�v��;iI���lxp�4Y�<}��Ns7�����u���N-�4�'knĬl�t��	g4;k��ٺz�����qPŰ��	�	FM*,�Tk�nY�F��a����>�o�p�F������,�F*ja-�ICJ�TDF�)ȡ�3�)�fX;����(�=�!�ܢ �M+�at�U5ڒ"��j-��� ��>�2��V�����S�v�6��c?�QW�Ęe'{ә:�؈`B�4tg�e��o�������OZ?A5]�W.s�A�-?�鋚^���oo���6���X)ٿ�r�o��~Q� ~Z��JH�:���>}������1�11w lni�z'}�)"���`��K��_��(�'a9)^�Sk7�r���#O�%K�X����k�[O�zt��xd뵹,��R���E_��ʲ�V^����`���B�����[�͉w.s$Qq�n|�Mb����0�ip�MHP`s<�
��n������ވ��n#>+L�;T�k5;��]��Q�,����5�+KH0������X<hm�J�,��j�NN[�r��N���Xd���-λ�>ZżWĉ��Yץ�ɝ�pL���GvE)z�G�H�:FGm����	!�E��LV���D:��Pf.�v@�|R�d�^�8
'�u9���Fĝ��?۔N�	)��L0�%֙t�-�`�uםc�ٱpdN��և�3��0vP��0�u��G!/�0����턝fA!%��M���/�7��
��&	)10���U[�E����ȗW2s8ɢ�r�����e8�%�b�cb���/�j��S�f)�����ȝ�X#�;9�g"bfe��T��$�2�CZ�I�Q6�����!U^�&~����|�2�����=�pu9�����^o�L'}R��8�u�bN�q��)Ǿ=Т����'6^�z�MQrBJ�M����G�2&���\��h�������nrT�F����x�RGF��L�H���{��E9Z�t��W/�,̣_�L�ݺG�|���z���}E2p9K��x�D�/0WY�0֖f_�ݼ����4�&,6����VWw��o����y�>��:�{��foOY`�?�GƝi )�3��j�k��bEљ�p^��צ��on}�ǎ=FF�ƃ���6�@�TW��^��M�t���)�k�܁$�i{�̄m�ƒ�����o���3�%�}}xx���`�����/2qe�);)K�RW�W�Ia�5�����ja4��;�dg�g�ݒ|-���Gʆ�ė�Oߔ����>Rt(Yк�nM�Fx�ϴK�}�<6�����3������2���T�ښ�Q[9]oo�jMk�|�h}�H�V,�8���;4 `��x3_�h�#�v�~	�C<��+�x�/�`�HT�
�I�}�)!<ĩ7 �퇯�0����<!�T�L�L���r��>���wa����T�!�^��Rg8Uj� �v�v),�eK^!��J�c>�q���v]��S�9�a:U3��H�[w�c�h5S)^��yD�M��L�iRO]d���'�71L�n�bb^g�|g#�+��K�Ƿ��nM�-���S��U��k�:��mʚ�^g�#��w���f��Pu��}\���\�(6�����m��HV���y-@n b|K`���*�U�ſ������뛕ٜ��XUTP�{U[V.w��5�ijޣUY���5���j�m'g,�n��Cw��&���k�x~��X�@�DBr
��82\yh./�.�i5�,���:i�2�S�`X7�CJ�+B�	��F�w�V>�+`<�#^?�Z�����G��kϒ�%K�zc��1&��8��_i	�O��.�͍k����-Wr�ì�<wN��׏�����:������=DEEŭ��R��I4��x_f~Q!<f��r&�߂��HɅ�n��R��@���xS��T�p~�d���x��ym��AN<�c������Y����[�/Ķ���m�4J��@3''ը�{��� |/��������o��`�פ{�Mл��.⽥r��Z	Ks=n����↪Ι�P:n�t��@f���t�tJ՞ǢvoX�̽�Rb�/J�,J����F="�2h����v0�EQ�����ɖ[X]]%�}�*,+c2`��h�:<<����Y8:x�=������,�}[�d,��X6U�zk���+g7��R���lI	���-Wh۩p�ڠ�3�9���8e��S�\O:靈������ׯ��_k�p�?��&Y�T���T[�]�c��ӗ�r�Q�8��_�a�<瓯�D�x�ژ��ۮ������N^/?�<���!�.^U����I�d��p9���Q�G�%=dz���4)*#�����=��8;�R��	6��1~�}ޞ�7�N��@�a�g�ݑ�Qi��x�6=��ʜ��<�+k�ںמN��<��;c���t�r�k�]�>��COS�#�V�A�3*��^��GTW�5uʓ�4���>���y��q��a�uc����*����U{?��5,�f� ˰��Y)��y]�mͭ6�L,�֫o��f���Po�ff{����+<%�}:�9(4Y^ 1� �����NrW���%�}L�)�p��<6��{���ld�cݻS�ب~a�	���"����K��}�\Wee�Ur>ٟ��ՠ������G��;���k����\q�S�S����1�徬�0:�[\����*8�Il��I_�x��@rr�ǟmat���a<lV�D�d9��:ZU��s�F!�e=u������2A���_t���tM��B�K��dmfZf�J𸸸�ֳ�z���p�i^�����rW~w�u����f����z�z7h#��[�:?zw���j�s�61%�����1����u3K�2�����`�(Ɉ��>���/ż�o��ҿ��!2��)�-xd5AH���ʲ�0��Η<&��A���+�&o�'�zz$2�ǯ�}�v�q
�o�o��t֨No= 
��)�fШ)̣��X�j���
��W�1F����Bag���
E@�0�㢔��ѭ��15��̽��8e^x>�������킥Rv}9�����J�Tx����}��������	��-��ۙ�>�uW�k���n�c222ǦC�$
]��򚩆�V��%�z��̰|S��| �V��JAO�/����v�|Q�-��mx�2��ׄ �  ����I/�=��"�*_���@��,(
^|u{0��nP/�����v�x�2W�2���N(�4�R��[��p�┉�v��_�D9���I���{&!����<�K�'��`q0g�H���P{Z-��������`�(J@Df�T���ג���&&R���8��חӳ���@�Γ�D���R��������&S҃����(�hN������|�z���|v��k&mI'W�JS,p�P�Љ��_�:o=�ٵ�E%N���n�����o<ކ�"�[�Cmm�QF�վ�@" ������g��Tg�blc�i�gWZH����w�efN������/ Ұ��QϾ�����O/ӎ��l�p�_OT}��f��ogI|�	1f�t���~�k�㭤��(�xyyid��abq����9��yg�>��o&v�\�;-�zM��Ʊ
�&��`7�=ʑ�k"�>��#��emJ���r��y޸ ������x��d^��.���ԠCC��D��[�Jy#�1{{fc/pZ�_2�dH}@w۹� `d�������l�Qx�Gr�3j�R!�.�c��k^CIm���T�ݪ��%!�M���x�55c��e��:h��-�L��Vq0�kj6 ��d�Hc$���w��ٰ��d1�atk��錡u�{	I�i� ��Gg>�rNbB
sdB�:�w�IU^�^̪]��������;��r#�c�*��(��k�7?��Hd/�F��?�dQQ�g}}�$��'1�"2��$�����mZz� )��h�4�����1ǳ�v�A�@����\����:�-���.�)�g��ƷNh��u樏�Axv��G�x���d��
��/�)��&Cp>.ܴ���[�]G�Ϳl\8�E~637��:v�܁�M@������}FzU��h�Y��s�r� #<4Ku���!�}[�����ǳ�dx��o�B��M�˷L��o�Re��m���󵒴:-;WV�O�A��Y�߿���=�T�IT�� �[�61��H�7�����G�z}�N��#�������]�♡�����@>�W )�I'�����mB�� �̟Q�t�����ȎL���uBp��J��0���+���։Ir��d����ޒ���	fJ��B�l�w������<��bƵ[�"�~i(E�c���f׸�&��彩�o�\k�f6,��m�������KXR��7#S�V��S5������&!����FTB�D���߄�K~e�䥚��� #��Q�&XD���ŭa�ߠU)5�fB���9��w�Sf"_�{�n��$w=���,��n1��"	�$3J'�;k�� �\��/�ˈ_�������C&3}���ė�Ny>��胸H=`թ5����V*�������R6���&�p�:G�J��y���Cӹ�tx�,?�̧_�R� �̷A%�m�]�[�_�K3�Z�M;9�`��[BK��Z�\ h�?��nw�Ս?M���������qSN�2>�症&~3�	�Ii��t��
���^}.A�AL��X �| ��L�L��YD�H!��~�]�"0d��nBÖYЄ��@� 9|s!3/��s��p!F&n�k�*�0�f�O����\#�1�)��H�;J�t-sr�_�,�����<��xu5�D��:G�񊓎��<�]�u��W��Y����m9)���:.����e�Z��Q���Y�$��6�oڌ+#�mY�m9�o�:!8\/s����fD�~N��Kf�|g�a��-�%��YC�-�}�}�M��9��]�K�KԩV�U���E��R��,9�ɬ2�%��kK���?L��mh�s��ws���D�6'_�)�ǧV�hbhX��XdбK	Y@���S��m~]��O�#�ߔPCbnt֢)p��*)��4/}_y�&�Dk�z\ot�~VL���5x�V�D���
{;�u���-�l��j:B�Q�R��M���x�ڨ}�y�66[��ίy�U|�hW˟^���������9�%�>H�2N,���K--��Uf����)ٜ}���
2/nk����ϗ4����#�:T�6U?��F
g�զu���w<<��.��G^������;�	0�g����e{�pSX����,���8�\%�{J�l�e�9_ϊ[GB����D^�!�"HL��7W'Gn`.Xi�O5�0���'�0�v�����ĔXz�j�x�j��ƄԶ��;�;�8M�C��`�[�iz�4�5@n��3�$i��O�<Cc�j�4��+�����!�,E[����_��F�aN�+����
m��]WN��A����F3ٙ��.��D��C�.�$d��1�3>Md0����Н�4�*|7��7-�?�9dt���{;'����ᑇ��0'	��Gf�U��Wc+h��$�n?h E�E3�f	Sjw.��$��a}m�J�� h@�g����6t������d�������9G���_�[Tul�c����KK�WX�F�!^�}򏢅�6�/�2���
����>N�[������{z��2K���K\;h�4�7jL�E�C�x.�4Ê�kA �zq��f�\J/JB}\ʜa�@O��,�1�%`扲4�%��F_J�G�Z��z_Z��0{�}�\�]Z�^k9z����an���\�#����c��Qh���A�W�U�+����ag�Ȩ��Dh�9|_
��x�S
��@�����'������ɫ��(���{?7�>�G���i�=����-NJ\�&���vLȪ7��f��5�
L���}�ttw��B�K���V4�������� �0n����e#t��	��u���o�8\$���(�^���ѻ�DbJ8&�Ț�/vN�#l�e�����Tq��j�޲�>�Eښ�F�>/U:}�g�&1���m��g�4�_������²�����3����F�&����齑�௉-�X���9N`��;O��Lk����Xx�[3��ǹ�;��)s����4h�jR_����/��'"lU����2�M�5"�M��.5(]��-]*���mqLE{L���H��cH����A����0�/;ny�c��ZA�[R����S@���8{머�-|0,8$���%�� � �[pww�w
�$@p��C�N��$4s+��~3��̚�X�Zun�{�w������w�2_���R�ܧ.��k�u�%�C�]!�Jku鵷q�O/&��UAT�I&e���t�{�FjX��o�{�U��^�5#͏Ņ�,�6��:�괶�e��%͏��dX�x�?��*���z�ѐB�C�[i���|(�ߢ�>��x�(�F�cvF��y3�cS���'��ED�i<�8�φ��GBy%�L��u��u��22a4����j�C�Jbh��dG�R��!�BDD�	������3��WsRr2Gӻ�ؘ&
�^�>�&������@A�/U��bA��P=���e�u�o�j�n��C�}Waca�|C�Yn��9�\װo�70�ƶ�2��g�jyY�H�E�`�R�*aq�[�Ee��|�dˀ!���>�F� ud�A��@[b]_�m{�e3�'�c��'j��ʦכ��D���E�������=����{]����x;sYV�ᭃj�-v� ̱�o&/	W���TW��������D�WO��j�Լ.DH%��u��1����s���f�ZG�s@W�WQKS�>*��dȕ��F��ɠYz���� �@r׏6��"6˲�&R3|��\����xh�"� ��K�E�k�k�}�Q�'H|�t�W~X@��������z��u��D�<�[��*oA��{�L+�����z�kp�_�gu��c�c]��%߇�D���ҧc#Ӓre��b\*Tu5�6�t�z'�pwp&%�6�R����޽r<�
�˷���
�/�&��/����ʭ��M�qH�\�s7/o:%A����s$JPU*;�����1';;�g�n��[�Q���C����m�%��9O�����P��^<R�a���H\�>Y���Ie�8)���;2*��E�U�'���{��H�[w���a�:���iAW/R�FO��{��鲒76�]>�4�Ś�� H�<�<��-ǝ��1[�9����f�v�@{���B^Y5��ܚό�o�Ն�]�# (d3��������,�qf�F�QH5������K;R��&j����E��r&/ȕۥ�5/9�Z�閃+�������I���e��B�U0D���X0G�h���Lʥ�3��[�/�r�}ѕ�4�j��zp�n	,�js;8���./�	VD��ڳ����5,�@����v�=�+"?�-�0�5������{�
��Z��Ob��ͻ�Ļ6�2�s����[m����i�e	v1�?�'r�qŏQ?��!�-�b��UԪ7 ���}����V(��)��l��û�c�w���3w�Hwd�D=�2���<���$���l~�|����ꝻKY��s��_E5vO [-�뭗�Ԥ�\�����C���/�-
�p��_$s�j{��8���{vy)��L!wEQX�h�|�yAC���R3mWW��Kdd�:�
B����aDO0��!�P(��<�����ͣ������\]Q�����ʈ�8}$���N0޵ٞ��9&�>�����k��۸����bحwd:u�Z��9��/�}�/�=)/
����*}(߱�lF�� *��.؄+�8&�r/�)�-�����֓��z>���0Jc^sc��ҥ��1jߵK�Bְ��],�,���Ӊ�gK�������5z�/y9k�Aܱ|\��"a�R,ӣX�0�����
����xc�>��E��/'A �&���g�*��!ŝ��eˠO�+�b=�1�;�
v�:�>Ȧ/`V�w�����ۂ�q�ct�.f�I���R<�ċ��Gq�jv�[\7f(���wk�<!$n3j�|&�I�ճK�j����/�b�|�:c��P�v7]�W�s%n)9�Yl�7'��������O�҃|��A�=��=?���s `QA������*�.2��KztU����NԄ�J�N$�Y>�Ŵ�1�;�<D�&�^A�8~@�ڊ���T6�W�!����	��)�*ھ�i�����!UWz�W��3�v��t�~e�Z}R)B^�ˈ����j�PΠψ��s��.��#$D������k/�˲����>�V�\JI�I���zo���QZ�*�?/�	��)Ǌx������N�� T�Y���M�/�4�tg����c��	���U��"�z_���(�6�5���;}R�gp�������O=E�نW�-����k�iK���xH���O�g��.ϻ�q3oo&'��w��l�!�}1v5��X�G��feϧE4L��L&���|��2q�:ױ�2�W<���ZM1�I��WR�������/^��=GG|�H� �qS:�(��:%�j�f�A���a#C>�RF_YgI�� �F�1I=w�^~c�wG9���L�PB"��=<����N�T�؛8�k�9�Z���
Dϓ�}p�3���M�c{Z�#�>���Z���z��9$���(�yt��u���mbzH�奨E�]ڽ{缕������\s>r84���k_�~ݕ�i�-�6�]�,�J�|D��[��oK�&����לf���]gZs>��~�N0�|��ɺn#���س+��}��� �C���q�4��?~��,7
eh�~�[ӬN���e69�*v���r@J��'N��p�EGҺd�I�i�v���n���eH��� ^��|AyuY5�h�r��r���#�����]u2@�tTy4h��D:!'{쬋3?�?����L?�dΚ9S&OG�����ع`Z���-,:�����gBc�����ϝ_2�D���ޗ������ٽ��"������^8�W"z�mP�48y4.��1tl�P7sV<q�H=	/U�(����і����0����㲐8m=S�ڵcW^�=��	Y��o�y=�t�%E}Fb��u���ռ�cѬ�+S�E�@��~��sǵ	%�yNx�w�Z��y	kBk:$dg��S�V��ɪ��@-W)���r5���ϵ1��U���-f83 t����Mp��V���o�J��wM���4�>No��f�k�7�pT̄;pO��s�"���z�Oݘe[���|�����d<iɅ�6��G� �}�g�������"��r��!C�@a;�^�(��/Q�g�cj93_��@qQ��$6��'��L�����e|D�g��~��Q������gG\��)���8�R��\}Ȧ��ȧP��Y�K���*[�S�?X�EAH���f��gr���7Z��,Y���A�� :�ȸ}��!Ý>���������f��6��.f7:IհF"�S����`��]/lmywβ���2qj ����ףb'B�v�OI_��W��u��J�Q�8o�@Q�:*�-@앦Bs�N���O��P<�l��fJoe���$�x2 ��={�6)~ �(�w�6���ό^e`XAH�,�
L�Xw�
.=�<{ �~;��$V7�]l���䤞W�E��R�C��i�W���H���V."�d訃]4܀0����!�̸������5�j\���-g��Ĝ���nA��%7��˝�#���ǽ���E89)�lٮ$���/��p��w��m�o����VO{�3}�o�����|� 	w.�c�[~��7(m���*��_�,
Ie�D$\9|N1�vR:�>i*<畹��n#�\\���~�%�� )x�`�����'�O�_��8~�(���_�����ς.�W0xG;DUy��.�{M:㚐/�x����P�q�*�@]�v��Εd�.���{�1+`����tJ��G8�0+H��e*\����g�֗�.�Ի��p����Z1R2Hғ��vR��:}��k�1�h����Uy�j��V���V�!��\j�ĥD�LdN��cJc����̔W���Q�d��s3�Ih*�(۾� ��]�]����%��{�zB��rڇ����?�G��L:��a}7�w#�=z��5O�IO�(��L���h����Q`[
S��N��[����K_E�Dq�b��V�2,D���ێ����	Ǌ��#��$6�QwQ�x�JuPЏ�L��� ���� �[ 7�]�LMx �x�(u��1+�G��k�B#uX��8_m�X��ʜ�������l4����N���siۭc���g>�}=o�;y����_|�5�8C�!��T��O���Z����`0S�&
����A������eP332�$ ���g���'@�'��e����d�|����A�F���?I��:�4L����B��m-:k.�f����m��CC��X��`nlbS&��~��C�6MɇFN<�ðo�#
��%���ק�tG�����:�ct����g'������OҽK�l[����p-��� �N
&xU���_��|b���gn��.�c���J�2<�4����}�bR�M����.?o����k��ҥ v�3�|pU\�L֍�#a�A��vP1���%��~_B�9�Y��;��
X�����!�ǂcS뉓�v��I�3�8P5#�%�`��.��/��Jr����1#.�f�����(�I��c����o��W��i�KYP�u�W[�6n9���H�:�x����Q��VE�X���%i����à�.M���ZE�!��d�mp�E��e`���ʢ����$m���xx�t��������O7��(� 
��g� ��J"z�8\r�\��pQ�������{EQU��t���X1Y�RjҞx���7'E�	"�2}w�c;i=w�=="^��F���c9�U�x�8�*,k_�V�&�u����oS���7���skXk��1OB��#�s��l_N����L�s�ڤ�e6�� [�N���b��m3r��p�zx��V��K���AW��5�` �6\�W� cs�^k{���rT�hٖ8[����=����!
{u��e6z} �;6t&��;w��`K[�	�*x�؂`9���Cv� MM}~)mZ��z,�l��N���-a6�N�Vn�L����ر\�(��×�:��L}��I�jS����z��Ý�+>ifX�<��Ȓ��z��2�4���a���Z?��Q�5�g�T�|sv��}}F禎�Fo_+�C�/`��Mȕ��)T,��X�~�"ݬ&&1�+6��A����ś?C>�����p5M� ��_!H�{N�\����	
N�5`�Qq
����0�ʞ�8�Y���8����| ՛�N�x�����J��m��9O9S�o���[c�R�Ī����!��CM/������v�1���%]_�[���Ⱥ $ܕ���6:�. �=���d��ov F2�#M����0=�qG�KG�Wd?�"4v,�0��mm���!��4��n�2թlP~%
�{젫���K��yW�
޷� ��������|k�@F�G%1�M�������r���?$25�N"���6��E/N��H�a����:�y	��>�nz�[�����f.c��r?;]|��Bc�li���ObI�jc}1��zh 
�	n���0��dɝ��2�,�<�=������W���NV����VFJ�Nǉ�x�|[����ыzq��z���K�e�=o�f_{���@Bf�}ӽ)��*u���Z��W�/���؄���	7Zfx�V�80 �����Ui�Լ<��K�8n\I�.�¦&-b8-����2�vC ��B���D=������$�J�	��EJĐR��"'k��2�~��R��l{�	V��`L�Z�uA�(��}D-NF�Q`?��� 8i����}�� ?���ڹ�+�����w�����2ݢ���1�� <mnCavv��V�r�f�^�$&��5^X@ʺ�3w4uL	 ���9��@���k��ȌI[����I4J�j��Ѓ�N�js�غ�JDgJ�n�o�k��X����v;(B��-s�����:jwY��7ZX;~��2��F�4sU`c!k [���F��X�'ϝ6{��N@n%����(�nXW��G1#����S�V���O1�����ɰd�l.�t$�ʲ��,�O� �{�e��2ʁS�HR�x�ǀ�ӂͫ�[JW��Y�a�:�Ĝ�_�b��E�~=8C���w�3��.�� ��	C!���LG��l������sxj{��	hߊK���MU]]]'��(LM�������}N�R�ϓ�/�&�� Zi����?72�'��
��@�� E���U��K�4>�=+e��w����\�lc\��2��僯'�Ϻ�1%u�L�u����D�?PQ����7\���˷��v5���nC���V�m̦��-(C��&$H�*���K��GwȖ�.�I���Q�ظ�� 4�ቊ�ho��oKt\��7�GN�|_�u�k 2:�f\Rٿ��{>�����
���4�M5��8����{E4`a$�4ʦ �⢿=���(���k㋅��2�S�q��m�u��i�|�����s��t�˫lNM��	���T��\{���k�R86B�t�q?:��Sp�K���e4u�7�bu>�g�\ە��׻�����:2��K�/ڕ�z���7U�L�_���	����>�G�hq`A���������p}ϻ2�,��|���}�ܰ9L^k.M������ӹ),,�I^Gܢ��F|ܵ���+v��+����x#�����w����{������:�'<�y�k�)�����y�F��8@�Fs��B�\�=1�Ş��h0!
�)�͸�i�-��t�'�Ae��V<��wl����`c��QC���ԣ?1�m2�
�{\(�������\.ٴ0>,{x�њ'�̾�j�g ���:|��"�N��ð���f���yg�-�Ae��[n��K�	����'[+$� "��p���"�3��S�8{���ݐ!��)���. !ʥ��˼�=��x�J�=<4��7���?�(p@�/�w��n~���_��/ώ�؊Y���h\�p7���Æ���Re���1�;�?@���%0�[���F���g�N�q篅(2:��T@ �+ﳊ���#��px�>xe���b6%�8�A�t.��2�>��bى�i���,1��g�ssT�?a�/������DO�1 �i��#�3�i&�����'�hH)R�����q�M�EI�M�}A���m"��剛7AB��Z'0Y�4~�Ջ���y:��ԍ��)�=�hY;��
�>sVazs�,�s����q�iW�*U�]�qVp��.u�~»�=��3@�ͺQ��[�	�*f:��l[�d	+`V���͊i�����{3?%�*�18���B�ЅwSo��[9�x�R>t�{�VgG���b�Pr�D���L�/m�<w�R���}�E�,�Z#�j'��TxGT#��+_�.�(��jZ����mwv+n�ъ��-�mm���8�]����Zo�0�Sަ�B][���үn��F�D�W�$�7���T�.�������X��p&��a�/� �u�p��ډ����He�=���qkE=��t�xv(��F�����O�	���������W��T4sW!rG���|�ߑ�~B�
��W~q{+:�̸E��ha4��Y�����K���� i@BHJ���b=���n���E{��Cs��M��8����k]Z733��ׅ�F�d���tZ&p�$�6���4�i?+�'�d��^���e�Ī�[�ͪ�ϟ���τ����_�퇨�Dw�R�:�l�g�Kޞ�?"�A��Q\�TtT꒕~�W2��ʏ��O�r��pd�F�� �e����0��c�����D'0-��YF.��/������: ��`H���������T�ކp���&�S_sgQ�ͨ]C�"f�sj|}L�䠫Ca�^�Z@�p��[��Y��=�M*&޸uʄ�|:��zj3�}�+:���/8޹�|�h���!(E�a^��c)W��k�{��:у����e ��u0o��3"����a�J8�yN`"�e9�lƫ��ص���Y�d�4���<�w=�%Uf�M�='��#!k�\�b�ʷ[��0<F��_I�.�t2�N ?���uW
��s�d�;�S�-=j�O����]���?軗�X��,�H��V�e0�D�����w��V�Y=|<���y�pжw� ��/Sj���l�<��n�� 5qe��֦��}��f�B��a��j�D,4#��5	����Ӹ����4!�W�,����K�_�'=R۫��)&ِ���U��	��*�hU�Z��C�A.y]���b�������_�
��,.+KNI!����
{(�{rx��o��mm$N,-��\%^\�Y��$�fday�O)�Km����%�o�CT�ug4��}c����~"\���	횋普���fͨ���!�~�F�c�������k���b�J��wg�\����o�4!Tj�n�?�>�KE��ٸk-F���׏Z�N`ز���&Wܿ�Q�5cϹ;�p>9ֿa�/�!����k sEV�)Bz�3((�\:IpGVH�:3<#Pf�m�m-�:iQ���h�:3���U����u!�p���yb$^��w���v�t(0[�aJ\Rr8􀴞}iP��u�J��ցaF�po����0����dk��
�V��x�p?����"�T�k�:ղҭj�s���Y��Ž�Lu]����F�4������ִ�Lq @m��pӶJ+���S�lNj_�]�v�sP3����`��ىA]ջ�Ʈ���sԷbA^�ݪHї}����o/�H����Ԑ����� W�u��z`� #(dwG'M6�2�T]
*ȁ��f%z���i��R��ׅε7޼�y�h��Z�����ݫor|�)ӓ��$�߅���1��R1Ǟ=�n2+�z�Ђ|���/��Uբ�/�gM� �Y@�� ?x���2<<\m܇=���N*�$���O�$vW+|>��}��w�y}[]�9�8T�ɼc�'��J�psa;�N�e�.��8ve!���(��xQN���������ώ6P,6aY����'�sB�y��lSř܀�r���r�2�K%=��N�Q�Z+S%D�ͻ�d�f8{����m�k�֏�����HV�X����ڕ����X�����(��i%�q��m|�0Z��N8��+/57�����n��L�3g�-׉�4s�2D���܉b���yJp�t�s?I�/�2�kX{  Of��]A@1�G�b�E8Y��q�zӝ>�0����/��[��[�&6aYZ@�Ƒ0��se�浭	|О%��?��p��[I����x�Nz8)����wbBv{��@.��U�k\�E�W�<��l���
��g��bJ��%�H�Vy*�L g�t���̼��}��(�mB���؊/\9������^��Vm*�{L$�۬H`����f�e��Ý)��Q*%6�A����K TA�&�.��>p!���~�n4Xa�=�+g�ბ��=@��KS�ə�pss���dB��[Z����@���f��X����j�K;K[���G!�***T���f�QR�R\��ccq��EYB�_�J�)(C�8Y��Su���"R����H��p��y��������n�GX�&�'����t*CL(-�z
�~rx�t�"���T�x�A2�	I誻G�+�G�U����MK1�FN�7Q�G2�ڊ�Eԉ��� L�'f��|�ۛ�R�U�O�tJM�G�m�Ƶ��>�C��N�`}����Q#(��H���.��(���7�J���Jk�ɝ>(o�F�2O1�TҊg>��m:u4���nV1kX@�͕ݠK-(�g�SfF>k=��qm{ꤼܺۺ�YS�v��_[��-��x~��{ɕ��c��G�q�����p����4� ߮~d��T�y����"�
�q,�L7տ����h`o�m?_��+tX�����"Z�cӘ��V���>��oD+t���W��=�qs��e�"��V��Ƒ�7��L��_��� \����5	s�nj=����y䰧�4?�?q�M��2*C����R�$�u\�(|L���X�\a�
a:���:}0���16fq�H�7�f��edc57���f���677o��{*��z��M���imޗ�GЂ�&-++���Z5��T|����JA4p#ǥ���Y����U!�Q=f�~.��v��Ȼ:�7h��߭�,~l�߿�Iq�7�*".l�G�EOŲ���ѡB���Y������%KjdG^�r�C?�4���N�J	7�|	)bnVx1�à7)�Q��g�咢E郜��،�ɂgTS�X�i�i�������A�3�{��P`�F:lV`��	
�o���u��1��p�B��3s���^ ?��:4����[���=0��?�/�����D��R�P�t�Et�9`Ҡ$%�D��E����J��<Z1m s�˃��Lxt���e�e��[~�L�Jg�0�-}D��2���V����Fa��+��J]���GV�ָ�<&���!|SS���x"Ʌ�\���k�; `#�x��4���̫E�Ǿ1`Y�|�C �c�NY��xM�I��]�����H��7Q;���|5��28n[��`?�˨�R�7Yrn���EU*���X���e�H��u��!�-���Z�3`�$���KJ8�/2����9@~l�m��y�e
{N,.�p�J
�*��̕��q,��BHX�9�\�
�BM6�|��Ś�U���is?i��|�ҥ�NF4$tzv���Q�+�4�t&]jam��+'CW^�=9SF���j6%����rBz���f�3	Fj%��� �syl�,�(��9���`�J�f�n:<7Rtu�a�p��,ln�C�~�n
< Z��#�$L�g�5+< ^��7 d�w�qqC~�:�9K����"���]���Wf��wh�]�Њ�74���ػ�R�������s�&�S5�`��vsg����t�zm-]_�k�/�����sړ1��7I�tG�zّ2E���~`�k�]�肄2�^�SF��̄�S��3v3ZhQ�1�����CÍIt�^����K�$�(����� '�DB%eH}�Z@AJ��<M�~-�˦6�����S��<0υC�r>|��=��la�
���5_hܶ:���ay��l<g�[Z��nZj�X��u�3?��(��q�53�EB�`l�R���B�4T.)--(.~� ��|hC*@E��W���*r�s��������'��>)�^����R6�ƍ�2#���A�#""�_�?�(3�|���,k%ϴ)�N�sA��"�M��Ku��e_5[>'�fЕv�vOΩ���,a%k~s�Fﵒ�w.k�f;�\W���&Y�u��s[�p��
'I��X @Lkn��`N���p�|�y_Eq+qsY����GK�����=�^lNӉ<L�&�7m�9cc����2e��r����hK"���;<���Z]�U���I�v��
>�Ó��_��3����fT���L��"@Ycу^�Qp'(ma�̗Xҫ�����U���EZ�UIa�ikl�]��9����Us�(��aRy��<��$�R�@c��4�9&�H�k����  ��QW�6��ɣoF��ee�y�}Et����yފ���w���dq2��X��6�Th�o��y床_C�kؾ��OCxp0?�=`�����2<�ZmpЭI<�����|v�)��o���g��T�e�d���>��uV}���xl@���Zv�y�ͳ4����0����f���>vXAy�"7�����j��aU�fqQ6g�I�����1��6`\\r����)))ң�Z���GK-���x�H����a�|[�p�8mn��0�G�j*�>G��g���ztW��5���G��?�a �X��8�`��ƛ��Bߤ8�j����:<{���f�v�9oc�ڝɁ��pB�{��^C�L�:�a���!4}x�x�2���;�t3|9ܩ��1�t��0�k��nk����Q8���ͷ�H�T%���3�.<�)����}�Dh��-�8�xI�g��'�%��k㋄�����F/4y� >0�r���J�t!	,���q�A���e��YY	�ج���8�+~��e(�����;a�!.3���1�7|����/)��B�1�c���˙�`C�)�cs�Tq�y��z)��6�;����uʸ�4*m��eI6�q��}.7ߤ���:�p'�ܫ��)+�KI6n9#��BpUJo��G[�0oדwDv��l8���y�䄖�$�벡�J�0꼇A13���NV�3�Z�W'O�;���S�9����������'�D4�)9�	&����?Kp�
â��6��	�Pg��_m����ׯ��)�<�<]��KM8���*Gc���zEL(���6=�D�µs��]�|�Jv7:��_[7bT��J�̓����o�!j�VG��ig��\0-*6$��(���{���o��2�Ww�!pw$6a�4bns����h�D?�$��X֗E�,=���-*�:�`�'ͬ�a���J;�D	��w��p��y"�3=�	�B:�Y�K��ܮ筺�@{ɔݠ���޸�~��ޥ�y�l���y�ԟua B*z:�V�B�v��s#o,���I4��11J���ά�O4=�X֤�a�'٬d�43��8"��Ѩ�8�^`�o��	/��z3OML����<��r�0L�1�4��_{������<s��
���]w7�c�����f+������/é�?w�쨃�Ш�D�%�����m5��Ai~�~�Y��6�����N~��66e9^Ĕ��Y �o��g*h{3H���[i�	muzo&���Lb<q
�@�X=�����Ԗ�7<��"(�!�E$F���><<<���x��9�夨)�Iplj{~�Z�3\Z-�q���)rg{r�J*�~���l~�͗��Z���f�&I4�h�ۉ��������g_������9�6:�b��M��I��%w$|��
��|"ƌ"֫�q7�3I�
֖�)dRB�m�L���Y;�<����	�墔H��Դ������Oĳ�ێZ�ߨBv[&L�n�����݃NJ�K6w�?��l��m��mی��zX�*6������1���N�~��y���떼��X�+��F�sJ.{�E��܄��^mQ�H���"~�W;�6��.Y�s')����V����c�)ȿ]:-�Ïb��6�>�`1f�?�W����`"�rF�`��M�z�LB�����ϳi�ZAC�~u��g0�@6M&������RE��]+E���XCk�]J'R⚽7�K��*��zX6^�1 <�m������d��7�����"���f~�O.=�!���WK�{�*Lz�-�ƳXD%ϵ��Ϟ�[����b���78��}�\�YX����lc!4z�Ŀ��z'BaF�ns��'&[���X}�Ƨ���q��pq!!��]�w����>�yHB�����oUF�i�OG�?�~*J�#Z񤠣�;��N�	� x��w���B9*�RAQq��;22���V�K�Ա����W��Tz�Z��)������kff��˗=%}��(kǳ�w�BF�yX��3Vq+����N����wː����%bQY㯵�q�x4yЧ��$̀:��L��A�F2��ª�fv��7M�����_6���>+"'Z��_5(���ቑg\""w�ڗ{Κ��H~�a~r�/�P^�(�]�e�	�S[.���Ӽ�l���ƫ�E{�+�b줊�n)4
e�@�ݤ=>I�T�ʸ���ި改2U7�`ϳ�"c�~�ȳ<zOܰ�a;t�,/QG�$��f LH�~�S��i�Ĥ�2�;�������Z�NM�		����A�`���=V�%��c��9���"|��B�&p�9΋��
�h;�9�W�SxK�+�O��IN����_�NŦ{�O�!���^Q]�ǲ}[������Zc)���ؑ�����^��}�.cn~3��xs��=�Ƀ�R�8���*G�e�H�^��$��H��a��It,!B6���W��-B��|p�; �����I+��"�v��L�/�;T54q\H��s��(c؜'�''��%��B�y_�NT$Kp���prq��Y|�ln�+()�sh�dW��N!"��:k,��|m����D���4�;��nu�����l���_썀,Db��L'��w����u5V��17"�Nk@�$��C������+9��T�����C����AL���cjw ����1J�Ef����~�_x{=ݞb xf���a��C7L��t��:nT�t1��o�4�-u��NE�β�ϖ��T��
eDblX��I
*F������h%���sG�snb)3ssS3��?��FA���7��٪��O�6G��[�8�a�w������<~!O=���
xu�������(��N��u�}6[�Y�V^L���k�\��h�?>���Pr<������a�x9�ߛa������e;���Ӏ��F�^��;��Qy�y�*
��@@����.��Z|�/�S���|����*���XR3o�n�$-=eY�'m���Dtߑ�r9���C�ڐP�?�H��F��߇@�ۼA9׋Σ�tt2�@�HQ�x99δ����i��ᏸtͼ��o%�)���.��md�Ç��2uG\�X���u(� P����Y��H�?}���K��<�b6^j���=�U��/Z���I6���v�6]�X�P]x-��l�j�1�ԫ+OXJqjh(���=!�Q�dum-͸�����	�hŧef&��["�#z�*k0Zf��:�� �w?ȁ�h��M"���ˡ1����]��?i�fo����m�n.u3���ƃw���<�ξ�5�<�f�����q
t�vv#�aU^��(UU�{���7w�+�X�'t�)9����rh�"��g �}���4�T��~�v��B���
�Y��j�i�ǯ�����;F9	�X����&���7�����C�hqQ�E}�Jㅄ��c�,F��~6xҙ��w?2�WM]=n �����>ǲ����\�0��IKK�%����5y�I芌��3a���Mh�<���q���䁎���>N�v�ebXYZ'��1�f����dz�.[��[.��~ͻY�P/��/���Oϫ.�_?Ԩ2�<X�w|%s�{�f� ������d�����T��xLoۛ���<L
:|��ݷDN�Ƈ�ܝ�# �S���zuM���� ��l��vG���r6����7� ��=絲�4 -��K-�:}�w��	�wj-�EJ���J��}��Bki~�xH�O�ž�Ԉ�� �ܼ���X����U`,��D�1�)�a��_� �P�o?�U�.�)�ȘN[d�!E2l[5ă���� �M���pr�̔��H�o3����[vB��5V�{۟�C.���0��2qq�Y������z��q
��A�
?�r�"�剗uJK���xa��a���j�:�3��z�	`H"��s�r@��~ǫ|��=*D�=�^yJ���o�	����Py�Fb�+�_;{v}:�#[�ɰ* FZdrp�S[��#�Rllx\K�W�D�1�%V!s7������/Q��3��F3���4��+�bn7���(�L}�@V)N�n�'�Jr�4��x`����i���}?U� ���
Rx��}��~�w?A��;X�O�@�$������F�?8��U+)��#H��l�]�mϑ|���?�C�MqzwՕ���3�b?��.H�tq��ovϏ�[/�Bh	tg����!g�܃�Cd������y{q�����Q��kx̜o����R�I
#�����?÷x�b��kQΟ�M|4��u�Y5�ʱǴ�N)�k���o�tS���&���"�H>j��u����[�C��*�d� ��T���O	Eť����x~2D8��m�N���4���!B�nY�s�{\��9)��i�gЍ�c���L�!������S=���w�!�r�nbK^/���J�ўaS�,��/���Y�ew����������pDVz�d5��� 	���1�6Ы�,绰7�D�Ĵ�s�4��-�>w����+/�Y�7K�/���
3!������� J��o�&��M��íi�ɔ�˰��W�6^�}0������/�r�w�&/ӓ]�S���.�u�=��vG��yǎ�G��xS��)��vsN�$��K�_�'�􈷭~�n�1�;a�˝�V���B�z�r�]s����Vu�&&&e�b�� �+��+���+�486_ r��~� �7p1�;��������sj��=X��
�iv����j���A�XU4��[��jg����M���ѧ�% �~
3į�
�M}!��C��|5���1�r��c�T"���\$Ҵ��zbB���Q�8�������7e��`����W���=o�.t9�i9�o��1�E��5�Nn�$��e#��9�V���"�����u���U�9�.���B��n#��%Z8q�����?)N���r��b"����Oe���|�1���v|�ŘwѶ7�Nb����i����%��6�j�v\��}U7����=����b�^����ؤ�s����"�1P�G��E��q��',.@T�'_�ݽ=��8G7Yp:�8V�;��s�Җ�.Y~�N�X�h�-��j_t�ǌh��8����?�9%��	��_m�~�&�$�8j�	U@E�Eԙ�ౝ�"��rY�H���}� ��eL^,�W�tq��P ##͌)<#<E�٤;x)�1:ն�W��o\Ԕ ��������%W�'d�Z3�w��ݗGw�U��|/M���);��"�;���V:���MK��`��Ϭ�<#�F���$*ب��^R�G��wI�ʅH簑aLR+j��v�~��|�W�G��s���^�r��k��+�߮�\��E�Ѡ�כ����t��#[�w
rY%�1`��r����oV���.b�D�o(�w���[L�6����٥#��,:p���Rd�M��e�kS�2}�Ŀu֫
�l
<n{-<S��0�A4֘��
D�y�Fš����@�ꗫ��wK'6�������Zv���f�9h$�K����Y�E�v{[P@JR��n�U����!�n	i�Ρ�[��r��!���}�~}�vߣ�qz33^׊�ֺ�i��7�KE��F��IG���p��E;�k+'ؚIA �1���=\��y� ���I_Ex���K�NW�ye���:P���w#	��u��嬓�fNx2~����8�,���3a>��U���y�|e�S` &�yN�[��r������}.�W���.s��*����#�/�Tm�?G#���ԗ���@?�%�{�ZP�~���p�>7���X�"-���7sN��r�'���+�<�^��>�dVl�fx����o�_�z֜z��Z���|��2�X5EDKE�I��	��o���+�,�,����˚��b���LN�HC��*dlݠ���E�D*�-
��L5�]�B�nAo��n�T~||Z~3%�J�R��7�l˗6�2� U>��Ð�r�
G��3��4�rR/yL�Gaوa��Kʂ]t��_�<Z̏	O�1�J��Ay�D B��pOA���$����κ�$'���ş��TQK�e�~��K��������ӗU���HY��v�J�$GS(h|hyש���@=�'^@]�F��ڳ?XLa�VґS�I�*��g��'������=<y��F�WS�*b��m	��x&^��U�:y6�#�+����ur//-�G�߮��/0˙1�{y��$�����Z�����A8� �H��Ar^����*�M �%(�S�k˭����I�a	�����������c}���G���ݪiw�V���	�
��K�Ǌ��}��=<=zz��KK�B��O��3���U�U;�K����v+�	��t}�H��v*"u�i�a^@��Y~�G1T0c5��R�w�M����7\
J�.;(Dw���4�EбJUr_��A���eB �ޙ^�K)I!m��3q�7��A8�u����Dux�)��÷W��C8D�rq\�9��rq{�����4\� �� �h猢G��7lJ�\�O�������ʤT�(�C�y2�@mj��� ��n/?W_-#����@��8��CGYq�w�o&�iy�?ۂ����y���r�n��\O�
sN�Rݯ:f:$Ș�a(��x��`�����ҶK�G�
��ly�����y5
�ܑ�4oJ!��^�K��e�,�{.?�8�`X���,�f��lV�W�K���u��;߻8��UP�g�LU������̡z��ʺt�	f�����m����⠐��FQQ�n�b�e;��Xn���h��|���u(�n�+��ow����g۷����EF����/?�:gz��U��._�p_e��������)4l�-��'��F�kry�a�U|��ϛ���M:�A���铉�[��e��c"���Ҧ3md�F���J�(p�@6�.�O?���~ϲӰ�Ji��.F'q�B�h��{^�2R��jz��ZSҼu�_���a�0��jh�P*�Fڰ�!�_ÇF����ݑ"6r�A�d��]<�H~ �kH�'�#�uz���N���L�̣�	�i�Ί�ڱ�@t[i��Q�	�۴��V�7�	:svc/�I~�zJi�9i��l��x,c�m=LH<�W�#j���(cա�) #�2CT�f�f�IY)s�2%�B���,�5ε8}�n����
A�������k����ݯC�&�~7W(��k�k��Mā���f���v-O��Aȁy����0�R_��<���J�+���<޵<;I?ߛ�����9j��_k��/b�"$5������-ʿ�晛�������^���1J�����B|�<�\���U��D��S<�hc0�����U{ά\yx1�	~�-��,gv�&���N�A�4�|Q"	)��\Hp�.�#�E�����6�zXF-׍
��\C<�^yŹ���G���@G��&���T]�����a�Q���KH�y08�_�~|6��3���iWߗj[�6`(�U�̗t�|�t�,Tܲ���E<���z���)!���O�f��z�B��ɉ���>KOj��׵ܐv/�0^��Eg�<�"te��:��ҭ�̔�Y�p=Y)���وdŕ�,�qƥ�:�nM��o�a۸8;��>�]Up���D1�h��́^Z
��-a�az�l#{��/5�I�ʇ)M ~������J��B�4@��J���%>>ALf�	|M?u��o�f�%5�D�<ȑ�����/���ʭާ>�;y�?OY����<���%���>�������:�1�^��w|f�)���<��O�?;�����WѼ��-G4lx]k��]U^⊅��o����,���U�����q#��wݪ��x�@k��EZ@��uM��q�/_WFj^&�i�M�^��*�23���&q���&E�bY}ԼBb�lX��M�T��+d>e�+�&t���֢O�g�������zm�f�~HuJ});i�:���r�Q�߉y�k�r
�ρܧM"�$���������$��|�|�>������`�ɒ
�W\���E�#��E�������3)�����u7z��F�S!{�j��c|�6Wj�QgJg��p���$��y��d�h����Cf��p�E���~�Ps�3��8@�E�sKDk�<8?{�73+�X �����roߢ�=t����V�(����V�~�.\4�x$>w:���[p����s�Lo���|�J�
R��"��{mu�s�ў��^���������.�xtv�m����w�ữp�p@������j�{76q�s��(���hQ�:�'���kAhC�.�⌦�?�Z���N�e�5*��{��s�X��5[��<��x�$�<��VUOM(�/�m'`j|M����;�V��\X�39�ᠬ����<�O���'���U�}�*�j�6�x�u
5�so��,W?bW��}��_��N�y����L���t�����=U�,3�̕�,ᖎ���[�P�~����1������b��˭���'�x����fٙ�:�n�jl�NQ���mmf�@�ݼ�m�2=�!�!4��IڨYLM:��c|�a�AK�+(\����4xH�[�>��|������"����Y�Ɖ}(��u�aQtp��bE�-hty���neYG\��UlI��R}{>9t�6���rj^���;��u�i�>2�ְJ'P��ʠCI���(_:��Ex�����C" lv�w��բj��i���dsz�z4w�N���ͥ�R -��DIr7��ˁ��
��'�����w�+ ����N�����&����_}����g��-xɜ��,����#��bȸa�\֒�H��S���7\�A�o*�����4O����s�;���)�>I�X�?D{4��1�\�XoDC�Nr�n=2Z��� ���d���:s,*��B�h�ݗ�� w*�9u�%�i�9���9��EyeKtg9�����CT�\�Vw����04�ѿ+��]��õ�CJ�L�U���DԒ��@Naؠ�a�a'���#�Y/d��u+Y� jPp������~�}%36�u�UL�
bZ�s"4��,,*KT�i:��|��<8��)�/_��Tph�,
��_*�?V�a�t��g�`������r?<u�ˆ�����U2{Y��<��?~E��Yg�����q��o�$9����U�]fXz��I��k�c��_>�e��L�wyWG<i��(��8�m�<>̻�%��M�������t��Z�Y���l��*���uA�b;�^�9�
��W%pk�N_���c�o�o���u�Lf����YI��|+�$�o4	]�^Y���풇�0���L�P��<��F��~K&�)��Y`�}��V����'�E*qrٚO��P��&�S��T�s�[��V�~����u��s�
_'�$1$b��/�P��y�\�y�7
s�5�b(7��M���G�� ,�Y�i�����I�ɶ��8j���˹����w�up��68�W��܏#������I��h0Z�s�['�|8������O?׃���cp2X9 Y��uv��rOh���½)(��./�/���"��_�T�Jd�"ɧ���A�)½�I>i���Yi�5�8U���$�c��(��.�ɷ(GڽO�'�<��gތ7A��WB-�P�H,��v��.%K\p��82b��W,������W0����ѱ&�%�4�k�X�`�I�X�J��y��%:�M�wY���ڐ2�l�PjI�`�ףb4޲�yetBs�w�/�u~+lG|Bu|37�Qp�,��PQ{�(Ț��l��078�-�����~�XX�j�ޥsYRf=�'�qU�V�������ϴyM��B��i�~��TF捒�;n���i�#~��t�~�;�G�zQZ֏v�8��L��%����׾[T�}g�T��"M�6Z�Xױc���ce�	�?mg�P/\�wo��F��gE�,
������\�
�O�sb����+�%��dk�
Ҿ{+̡XC�u�}�r	K�TX�9r��f���C���`���+$)��KO�m����!4������I�+������'7�Gi����t��)1L;	R�0��$3�bJZ�)�T�ݿ�P"c���os�]�1�k;9�5����������-]��
�k�����4R�F�f���.e=ē�qo���n��T!!*:�7M�/p�1ԝ�z6��H/����2��"K��6c�r(t�T��Vy�M����D�I���X�Xjϫy�pM�Y�k��C�:i�w*��Qmk�d=�����)�}��,�ï��d�a�8�/�oA�wِ�F|����h$����w���s�^L���݋���	-��,����Ͳ�	$&`������gBC��8��p�C�Դ��u:)�ˆ�x�z�^�O7���?���(f���Q�3J�j݄�?q���2�nlS����^���L: �Z�$Q�wG瘐0_S|�a��5S��^�_�J���ТM����cRR�-��7�864y�#u�����̤�>�,Oa2�����M����o�~&����w��A��	�(��휾݆�kx,�Q��#r����H��"�
wF�j�U���0o�����_C�	[�׮wCJT7�ȧ,��;��>����/e�5�K!q�Aԑ�}g�T�����jD1�
��p>��z|����8��R��Ms	��xVJ�9<���� o=��ەg��wɇ��_kZK�]��4��\ճ;,R;� �E�Ϩ�XW�)O�g��E��<q)Q��I�v�x���&��MTIH@@/$������ק`aQ���aw�u�(}�`X� �E�id�??�P�9�R�OI�
b�$��rgE$dVS��[N��Q�:�?to$�Չ;��R�P��9z�)mV���B�{���S|����z��#Ju�w��fhf�Nj�wޗ�r�5Zq�y���R��oo$k�����s
�Ev�f�.T+�n��~���}���f�r��ʒ�����ih)D�P�J�>ۆ�ޜ���� �R|�<��d�:,���}u�T&�[�&�,ν>s&��:�Hf/-Ʞ?�t���96A.p; i	S񭨬�IM-	{����.�BGG��u"w��ڮ2O%l�H�홧����t5O�J��)

�5��!��5[�Υ%��Cywߊ^��nƽ�r��D��5V�߾T%�O(�v����[�1̞�5�W}.���pQ�֑x�J�K�/TGk�O�k�臭4bx���A���te���>�.��xȤ�Wlsö��&k�[���D]��sK��Ս�52
����*١��[�wڲ�7J��A��,r
�ϟC�����j{hsDR__3�(T^����߿?���:!&����E���<c�?xΙ?��E �KV��v--c^I��{����m��EK]��f����#��0�֡OG�q��&(���t �R�@0]:��N��x	V��r���\H��������	�g�h��&�TϘ;�d�����w���o��������Ǣ6�\XK%U)�Ez�b��Cw�Q&t�%<�OӞ,y¿d{�?�^�||��%&�0��j�Ӛ�J�2�D�g��p2�FICӍ�ź̜�����#���Aʛ��j�`Kąd
o��I���,	�����2P�^l��9�˾1��i�8&�5�P��2t��q+���.U�_u4.��.U��P���s^Y�$�9��u8�\'�q͆#��N��/���]G�Ҥ�����3S)�3�nHM�c8X�'K�=}.zB=0�Y���|m4�%y�G��T���D�j�����z\i�������⃞�<��"�?�ōI��\67�cBzb� �������(3i����[�2����.㊏O�xmj�9x����y`��A�N]W���[���QA&��z���'&�����T	2{�����l2�t�*)��-��+�+�a����V���lߐ,���Tz�Ą+j�!�/g4d����4ʷsz��j��*�|�.�f�y�l�	SL�
�B�܄����N��]�`�~Y2E���U51Ʌ��"E''3��z�R�͛7^���7�>�Dނ�Ed?-83N]�>��x���TQ��`[�PWX�0���a��c��fs�4��XTZ��]c�قOc�q*)3����������В��kZ�nЁf��R�#Gԇ��!�-���ND{�����L����'JpO��@���G��W�H�(^&�6��V�T�m)���m�s#����㓕[
���0��K�ԙbP-/���4Z����N���e�R�#�P�4�oO��}qБ� %����}�9X�m$�V\IlllE#�����:��ML,�N���#q���z��2+��;�o�ξ}�\��x�$-���J��ч��OOW�d��0�/�V�_��5�nX'o����x�R'/��h�Vl3�q��}�\��A�f,�w�3�*�A	�R��Jv�r��̐�y���a6��dX�{{�oݎ)�5Nav�;8�(����`횣�v�"�e1���,���b]fe��^7�"T��oi+K62I7��6~��R�e�T�{x��ƶ�brkN+�����Y=�]�W�ҹ
?n[��86���Q�IqR�Ά�͘Na�G�gUfcO8�gX�՝��5�8Mn��P7W+�;n�P��Dj���Vk�c�`���!��"˷>��v�J?o⅐�t�Y�9�|q��˘9qH���\�޸Y���������U�R�@`��X�k]W��ԩ}xt�ϵ��U|��hE�Y(�'16}ҥ��n`��C#��v��rP �Q�򼵬�U��������;��f��Xb!���Y�!�F�q����n�m��0�ʍ7HKrU��f4_�2ăh��Daxm<��M��3����Խ�XP4�3��D�������-��R������ˆ��kΝ@u� ����qғ_lr{�&����4a ka�P��<�����-(|�n �Jl��#h[�ZJ�,u�f���a0������YEU|,��|O��;��r(�=�M���
�.�"�Q]��#K�G�I�s�{�<�����ݡ���`K��r	��٨,^3�_z��3���2��A(7��T�(�>sWy�3��~ 7���R��\'�u���ެHu���ֻf�%�q����m>��J�#���Y�����3����C��D� �ƭ5��;lB$��f�&LԌ&���U��ކ�/.77;�;��Sb�5`y�Te�[M�FsÚz�u��RI�m���X%su_ȝ�������+:l��ߐ�:���Kq>�Q��+��&O���As��g�ª!���F�T�Z��+�ïJ`�$�LQo_�6mA�$z���f	�m�쥣Wb;��׭�XoΞz�?��k�t����7
�ܭ_�<�U���6���w�����%6�$�b��˶7\Ն��;'uo�;I�����uhV.�ϒ��<)�Jjh$*(*�#:i��v尞�fAiA�?_��[4������ q���17������o�S��l�G_v�8h�`���Fj,*,	I����F�+~B>ɉ�u���uУo��U#��Q�X�e����X��JK�&%A�2ē�_�����=��F�Z>��gB��9.'hMvK*����l�r�ߩ��
NQL�;�	#	��MJ��[=�j�����vg���O�wjZ.T���^��S�⫛\&C��� I�I�V�0�4��C�Q�d{�=�{�]b�2����Ԡݱ$ŵXeO�x�V��0g��or���q�������������!�w%l"l/�"��ގ.�҄r�/�1�xgt�Z�-�	bn)�*��:������y$�L'�gM��C��BW�W7���f�ʙ"��/_��ML� h��ed��)*)]5@��sZ�^�}{�m�>"���y{�������?)�VTG��ѵ(��=>��[���G����T~��.d7��ܟ�����f욬�ixU�I�覊��ФL����aP�2���"��۔B��2Nv���M�M���p��;=c�5�7�-��"��H7�?��ڷ;�"Uy�dѰ�k�ęm��>��m������������*F��HA?\{Ӫ�z��`P��Qu�c��%����o�l=��iؾ>}��+q��������`�ҴT�Ӛ �W*��I��ʻ�\r�ֲP)b�u�HvǋӶ�f��՗�nWo�=��LDn.�!�*���5��2vt����Ў
�Ж��N��Pb[b
���mץ���������rB��� �F�Z�U�u��4��>=H����2�}����':�{�SE���qf�8���Cu��y-��^f����D�VVTx8�1�!���)������L�<8���B�fKj�0f���Bź.yh���� �r6f|����z�S�Ya,%Yٗ\بi�w~�o��~_���CȷU��V5���VS�I�pEu�e����l�P,�x���v��%�0�نW�S��F݌��J��6��:����ǵ�bcaͶ��aF�1�x��D��#�(����mj�\����4E�\��`;��7��٥?4���:�I�.��k�deLK:��j��zі��LI�c|�{QG��1��z���L|7 E�Ҫ�G�t��Ɲ���p~@%��\�rW��DN0 �^Jn&�uJZX��O��ﲼ��c��2�u���0���˼�N��@-��doo�%**s`@*��eY��a�1o3WqP=X��d0�׿���|��~������a���b��Hd�����,p�g�j$� �5%S1`pޘ~������*>i�� [�q��l��q#R~�E�/��
�ʳnTI�q ���Yw�|�W�ZĚ$�=��Ƣ�Rr}X��y_�eh��r;Z��|��"�1C/��m8��(����m	I����rn�a�� mzx�m4Xu��d��f|\�%r�/<	�/���1o�-��y����T�z۫ {|/р����v22=�ѰdS�J3�`?
~�v�,-��RbXZ�ʋ1������.�G�����S:5�S������Z����*��":5B���KJV��ZXX�%:�vؾB�y:�+�$�$�/�x<��m�o����B<xS�=|#��,��e�µ�3�p0��F���82�f�j��:)�
/��o�7�~���J��Klp+��>翀�%%�؝`���2�u������_ӂ(AMbU�����wԌ�	S��<	�-''�9�w׍ޅ"F��v���]Y� z�7�^gP�'*�%���.��1{�gKf[��{���k�%�߫e-�t��w_Qb{�a��XVjZB��,��ʥ�� ��܁.Z�����Q����jw���Q �oD2Mvf2���=n՛9�]�9���}��t���@!��LnffF�HJB"��O/*:���)==�$��P)Q8�\����ϞYX.̝����qzr���O��v*���%殬e7Fغ���)Z�X$oӳ,�~���n��v覧e��A@vs� �))�4:Xu�����Y��3�` �r�l���� 9��_g�e�H�3�����OD�4�+y%n��k3ǎ�{r	���E �SH~�:���F��#+�MD�d4���c�m�(��+��G`|�}?�["�ˤ8K���w�����%GQx�3DN�9�/z�c=�^�a;f��'����ri�D�LoUBN�J�q���r[^Mo��H���|�t'��O��gQ��&{�G�>�L���ͫVQ�r򭱞��⪩a����k8����Z�q/���2�Ȁ�����Dvܹ���lZ�U{���4Y2Α0,�{����~eC`5�����d`.��c���jm36����<��+:��-���X4�OS�N��U���K��=�w�<{es��홢99�7F��}����-P�b {'�Ts7��ęrhmbϩp��T]��!6�E7	8ވ�o�sT��(��H=�}C�e3E&����7��8Po1d�+ޝp/Ys}!3��������ڷ�5���t�:?���G�b���r��:��B,��,E��%-��|z��l=1h7,�Ý0�"l��E�����r����Y �`#��t/���@^��x֯����Ȳ�$Q9��T��Yx�H��� �A��v�/��Vm����v���}���wn�È��%O�q�V� ԟ�P}�Ъl�uLJC���,�A�(�D`{���L��aW���0j�^�1��`�~˷����P^�zN|�r��7�e4���:�d�0���u%����9����/�޻'s��nI�� Z��m���*:i]��%�9co]�p��P�m^J�0"�1j��oH`I��>�҉�XQ^y��7�|�~{�iqd
=.����AJ���Ze��fs@�6�6����f?�{��u��ƌ�p�}�pu�q��Z�12nad�k�Wm6��	�|F۵#���y[+�=�=.Ί㨾��L?ݩT����J(Ŕâ����}-���zĽ|�|X���������{��D��4���{iZ��R��˃�A����	�R���އos�����ɯ�Z9�XE`��!���K��:n��)�,��f�۫�C�2P�Ҽt_Y�]ݵ�0VC��4x^��=��^+GD�:2w���6E7@C����7��ǒ߃�,W����E���8�iEqYe393 F�������������*�=�2Y����Q�\�6[li~F���>=���oOf�A��.{݇~@�-�@+�V+t'�/>��a,���?T��	5$�Xƌ�V����%V�M��]��K��'�AA��L[�k�k8h_����x�[x:Lq'6����������ZX�R����G�d7#a��!���8��p�������9l�����R�֤�ڥ��l���uR�C��8�����2m-T����E��@q�������=]%������3yLY�(�Nyj𜹵���PrE�"�xx�c#w�J_>��9�ZR�N������8��ԙ�E���#l�0{5;/e��T�*Eʹ�K=6--��k�Z,�m�x�j]��V��s��Kgz�7oې���t4O�[#.
���e#'�X|*ʕ��D������ލZϒ�{�,���Z��cƒ�I��
�8$���v���-��$A[��O�N�6 %���d�T�x�T�R���ɇ���U�s�Cʥߴ�+7N���[�]�2�Rُ��C��v�9�I�
��םw�=�ê��W䃩��nǣH�\��-�3����}=\� .�n�QR��mB-��_��ɚ�Zd�2��Hf�0�������Z�k�$a�JG7
�?EΩ�v��;�0���}�O����Qaq�vr�!���KN����d�t�`�V�!A#�Q-��\�Yl��A�<����XL�6W�n&��bw�2a���Mz+�vP'o�X��"���Ҿ�FW
���/sCj�eo�5~�جCw���"ԴT����ܿ �b�K2�%5���/O��_�C!��΅L.�7�qhe���ď;��Äz��hB��V��	�5Z�%����nJ�44F�����N�wsS1`X(C�ãݙR���!#X�hH'rPQ�nOl'�Eƛ�����/la��_2�a���#��<��U�w�� �~wM5I�w2���Oѐp
QpP�T�<��q.ºGR��Q��+Z�Ԋ}�E�}����H��m�[oԩ<��ꡖM��me���^�̥�}dhԦ;a��\X���ZN���i�[3��	���#�Y���	���3�]ũM^��1�>������Eݕ\0�v��ײ�?�h�J�Ʋ)�B��	(9��Ѕ�*����Aq.��G4�'�6o�F����u���	��g+�;�P����������""���0TVw)��^=�@���y�K^����)��B��#(�<�w5�#����iGjە��a觫�<�΁q� �M��v�PE�������p4�"1$�.��؉�?7���Nf�`"V9�Y<�@�RY>.��m�P����< �kâ��~���bC�TY��}t���՛T�id$계<���>�L�����Ek7�A�������1#:��G�pog,j����"�Je���U�?Փiݹ�U�0
����cy�@��o!0��T���H�$�}��h�5^8�۷�kS-oX�,2|P?��+�t�S���G� �}�����#.^��ߢ���R�XkY�ih��2bU	���ʭ�6�fLD�,�v�
J��x����?��W�᫝�:/Hc�ۦ�a�wҶs}!��鱭��ҍ��s����M���+F�MK]�YH��b�̎I�^h_:
��hF���җϊ6+�r�r]=a����%�0���f/��ۺo����ڂ���������Rg��t�nCSI���u�kA8��I�:��;K'���wz�hlb��)�����6<>6���O�]��g��������{a������ISԤ]����L'j�h
E������V<U"N�����  Q�e��T�uyq���	��̸�e�oTe�$��t)�v���v�Y�ȹ�[&���R$zb}[Q?QG��N��RkEADgKӱ����ѻg{W�K�Q�u�Q���"{���!��3�~�.5��&���ƣi�n�k��bb��L�@��%�8�
��Mc��QչZ[�}��`�?.� HT��w�̛UeRq��z�=�ۺ5"W���'OT6CQ��KKW��%L�_[=���G�]�Z~`�`����X`�4�;>�z�������Ҿ����1dp�x�����L�6Ξ��אm�1j=C�8y�d��U)ĸ
��3ش��6�-s�֮�}�3{~}yɮ"��ߵ������!~�r�.6��~%�ku�n��(�^�c�����9A(�R��-`H?�UG��0$����oU��x����icX��#׭�I�ZN�����.,#@�	 7V��^Uq=��ޑ�&w��l��e���?�b�� ��<�&b���ʛ����*�"EGE wĳUVR�CQ������fѼXX�v���7�g�E��(n�e������'8[�F\G�*�3�KQ���%�Š�e|���!�z4+�)O�p��xaUM�X�]��D{$�S�ѕՓ�WOFL|'�3�t��������C��莘�.$;�:H�]�܎�m�����<![�MA�Τ�gj��7�N��1�s�b��ս��{
�����7@�F�1R��"�~+��;1+Fn���1*�f����p�v�[�u4# �3\�<R0�0y�a��d�O}y5��~����嵚����.�fa�������Y
[�/q�f��u�4��H~>(��9�j���*Da���,��IE=��Ǝ|���{"�4t.{� ��-�,t
���#�%��\�d����/)��q~����}�����
��`Ue��ug٠p�y�ܟ��n"#3[��֥7N&m8,)?݇��mg�ٜgy�&М���aH����������Qq�K&ſ�(x+w�'k�yT@!��fϼ�!E;�A"Q͊��jl	kl�P��3��4Y����k��Ew6]��BQ ��+q�OO������6*Jj_�˟�={lG/F�{��	���8.�Md��'M|���UP�U2���
�\#�	��%W��w��گ4��T��[t�����D�-~������R�ϒ��/!#S��_��tG��c(�qp��[�	+��}��y��d"��zϣ7{��/�c*�k��^ռ����ʑ��%pV�U��v��p�B�Dz����+���0y1���7O�os��%�K�=|�e�5�u��h�4-�J��a�d��cC~�d��g��}��a�k�鼷�6%+�<|�	>�0g������z��f�#��
y ���h�Z`q�0E�>
���s�\�5uQ�?���S����a3��d��J�"C�N��pk���������"�o=�j����Ӎ�w�~�B��κsIbI�` �d�) Hd�P�T�1b�0V4\�0T�[J��L�6:X��3z(Vc���E���H�JJ�}�M���nc?DCSpt��G4Dԓ����z�GL�A6��H�����1R���lp.d�����|)=����E�n��{T���R�x�{����A��ł��vN3���sOc�ԩ�W�靷q�l���ֿ��ʮ��q��u�j5��8�dv�]�@N���i��7�*�7V�H4I�-�r�DȊ���=5^��0�����<T��p&�#V��f��8`��X,k���d�6����5Z�T ^K:9>��s��~C1����ZU>�%e�w;%��c=C�$US���w��^��J'���;��tп���#��0��ccc�	숗#�_�c�-���ӧOe[㱉pQE�CҒ�J+��a�x"[���W�{�;v��G�ܑE�C@s�@q���1Q�n�!L��P��caaN��6�.���sb�a�Ӈ�rz����n ��jJ��hHh0��`��E�� ���LkR�~)F!��p��EL�ս��,;?����:>���yӽ�&�h� 18>�����N��Mv�'YH��j8LR�nWY�U{��i<���1d� D�j7뒗���,a�#.�3>���+`��9��L'7,9�D��z�2������,���c������d7E0r��:N��?4qΗ�5���D�D�8]�����[>����_��B%��5��	7�	�/���2'?�[�tR� d���� JqYfO��ng�tԳx�q-hX|=۪Zq)`�y��+V��kOz]�\LC�\���������xPֿ�5���Z-���;.��?V�r
#���;R�����qoŶ[��=����KLf�K?(�s����y����$_隇��C^@�'u�1���,�Mf�b��0����|	^N�� ����^�,ŐЖ?�3+��$�^�*U��渙�^Hk�]��q9;�F Bt�H+����4۰�YG	��X�p[O2�S����m�.�t�{m��b��?ã.��˾1���*�UJ����0ϧ���,�2�� ���3D� Rǯ!8��X�f.׋��iǴa7�������u�*z|�/�P�Tw˾}*��M|ƴ>IXي�l�"��z
��M�2�^	i�G���U�{�}���X(��e5m�����'��F��#s��3�e>���+��3��)u_V���W�R��*���@0<��
o8�v������oD gr�o#x�߄~�<!��NG���k|��w�xŐ�bkR�����5T{Aj�d�s�?�����Y����n��"��;��zO�-C��_�0�1�(������^�D�9�F�m���Os�"d_�g�����rE>���&�q!y���BW��觃��z-a�vC�;�@eK, "��4_kj��s¥�l�������6�<�gL�n�ߣs��Q+�A�\'���#��A�L��lb*����.CT��
eg|�3��|wrg`+us�Av��Z@9�{��1ji��Q�k��O�$l����V�ٯ�pʀ
��|
���	��{ec/ Jz����a(��D3ip�����a�Q���vS�clE�5���)����'ͬ�3�a�ܘ�X�JC��%1���)vf� ��&��~]����y�l�"){��K�Ck;}B��fހ,���\���y��l�DL�t��g�O���tl��@�F@��A�K���~$"�I�c��V7Qzv���ѥn�9K�Z4�¬	����XS�bu1ڱEJ�fK������������I�Å�%77����'�5�\Jg�z'�o���l�v��農�Y�\E�߈P���\�R[��*j��
�u��N���)�u\U�h��rb��dW=˩�>�W�z%$���^����y����/�AT��9�59�H��7�He��#B��=ܫ���CDF���M��{���|R������#mł�i?%�2A�e�r{��;N����繣֣ᢹyo�ӫ&���z��=�4s�:3�1�Y���㜚�q�j�H���)�I�b����HfÑ@�OK1uL^^����U���\�i�[���؏�x�p#��_���*A>�`����M�fԸ���� �YX���xU���1ـg�2???//�A�AA������qW��h�0���f����Oq��l�>늢U�Ht�k����Ʉ���V=�Ϻ�d-��Z�x�fc���阞�z�C55j��n�Ӏ�ĵM!M�K��$�Fe����ּ�[��Aw�.D��r��n��q��C��7���\��὘��T\��|�W���:M�G��V���w�&W�:�nD�ޯ�]W���f�m�j����^՚�:i��ω��=�X-��5?Sgcl(1��X^�N��.>��ͯk����������D\j��f�5x�3�#,OqQ��"���[L����X��*�!5�[v`�H�a��
��?��WpM,q�cMy��el�_��b���$Hx�$}�p>-�!}wOJ�aXRR�=dt���U�����8�ʨ����@ ����	��w'�[p����{pwww/��a��~ך^�=�|���Quέs�~d�}�Ѧ�����f��@Ƭ�%L�K�;tqU�Qw6������V8YT�wH����灩���!Cf�6E#�d>Ϳ[�w��a²Ju��;F�L�Re�=�>���BbHs���Q`m�Q� $=�V��TGV���0cr�)rV�#���9�K�w��h�,�xf��uZ�֥�}����#����˶������sZ�ظL������e���)�ە��Z'σ�2T��73�V��N��>
���ȵ�7$(ӵ�wZ��/&h��6���{�`
*� �����\]NB����X��K����T�)�Y�%�����1�<�i�xQ+�J�}l��(R����,���j���l�c.0��E�Q��<��f��F"�͜<�rz<�`.X�����S���Zt�|��[��Lϰ��u�6GO��O�C.r�0��"�P"u � �彠 ��إ���LrU�r�MN��V�J� �UC�a?�tg	�_��YӚ~[Y'���,��ϣ0�ξ������%S,��Șj�4>j�MM)�h�$�c���=�V�Dk��~E�E�������lF�^cZD�Ј�dw���ӱ+A��".yaW���#�MS!��-q�CW@�,R�ICL��z�˛��UP$&V1׋��4��,�]ӽ�M-�d��j&�q�#�D8C�c��,�����]�\N�����t��+X�5ůp�Ci����p�>h�.���6>~f���Z��@L�,\:�H�+C� ����9����� ��.���~��	3�"�kG�T���ַb]�ᶱa���+;����h��S�E4уؙL�}*Y:�O[��+��ɧ��Hp[ݗ�$���>{�2>;������ҫ׏��+�k�{����0�v��I_��l4$H
���'��5Κ�E���a`��U)UC͛霃�_��|6�J>���Z�[\�U���5�珘�l݇^�?"�I�yp�m��'��|��Zr�{��x~Y��)B+�������^/�R�����faP�`�>;f�+�U�9Qw���+_��3�wwT�ԟA�y�.�d�%�^?^��>��}�T.���.�Mx��E	����8g����m���;�K@���x�3�w��]l8C��~!����U}1�*�G~��n�~�k�Rr������t�w;�|���/$�7����$�f7T��Ma``��Z��n��!7.�$����Z1����]����q�Hߏ% $�$���iz�ނt&U�D@����2l���P'E11r/M��f�04NA@!-W�[6�._$⋮�E��b�_s�w�-����O �����(竀�&l�؋��ٜ�S��Hw=��ߩ���-�@�~z�9pS�`���q�''2dΊ�U� 1�}�1���)�u	�a/Fy�X�c!M!�mm�q�l��j$�aJKK�~-�{�7C� &3����:�%���
t)W���~E��]�@�P��a���	OS�<����%�淥��miF�c�����~P2*?S\a_7k��K՗�C�(8�&���#YB���;�K��_����5AVh�.�FU�?W �
SZ-�������mB�8 ��C� �L�������G�zzB�˸��P�h��P�_V��1���hl����&E��X�\t��:�-@,�(���T�r��I]Ҋ��S��t�����eƈ�h:�ǔ�+�8㜰R&Փ��][?'�����W�wC��xrq��������&}#ܡ���g`�y�U�����--8FJr�Un\ܿ㖪��:Q�x�Ʋlw{��%��b�%�5˛W���2h}r�l|Ӎ�MQ�=�]������I��yY�J�l������[������ߞ�"�����Y��;�,V�������jXb�x��Lw��?\H#�+ַMԁbH|�7+�y_v��!���F�Ӏy�+:&�Fk�:��}x|W�'���y6���ۭ���ɬt���(�Se����`-C��%�2�+����?���E����p����]���YCj�q �q��xA!Q���X���2��iE$;�9�v�z�HLCe�"-G?Os����GX{1U�IVQNt�y�8�F�{ӟs�<֔���m�1Cym��!o�>�ݜΛ0���<�^�|�����o�-,���q>:����kW�'J>o?"pl����2��sG�B!j��דV����%�f�&��q4`���Q��#.��0Ь|��(\f%��aW�s�?����\�;l�~S{�y��)���jl+z���<_r�*�D#V�$l����P�x��h��R.xp���i�;|�G����O����=��s������j�S���ЫJ/�Ԉ�@)9V3U�=�/ΈH+�1g7�m�7"���c쳛e�ж��E��1�X`��鶚K-?;�����i�&M��pX���"-gIqF]嚵���u�y�?Q\`��X�j6u�?�Q;A��F>��P�eb��|�E�|>���m��S^�vj=��u��0��h�H27�'���2����r� Q"����ve�\�h����-ؑ�7���
V�^-�&�K�巶��BR�l&����������r�	kb�#k����3���x���6b�k�Ξ�n?���A���Ϸ��t����#C��#1qpR��n�>�wa��o������ȏY�W�ጕ��[�]���can4�{����'-������*��҂��踲��t����s�;-2�:lXzB�V���bP�H����[u�a�׏�g�	��z�0�����a ���0Pe�������f=�l��4�^%�r$�p|��!�7�
q�����ǔ��&42z1�a�gN2Β�%ʹU���AO�D���S�0w�~$�f���s)���4۩Ef�����أۋ��d�9��^$�Pȕ��YD�;�]�W�kAz`���0��Қ^��CL m5h �V����F�l�(h-U#g�,bGV<ݐؕbeR7k#H��@ZBQ�b����1 m��Ll�6Qx�Ѕ?��g����7f�:9E{�$���ێ�}�y�&�B�"��M��zL�_�Q�bL(}�9�͌=��\3�O2��m��᜻	��Z���O������ S24�^�%���[l�J7"/cy�XN,�`�қ�n7��CҜk|8��?�!<�OGtP���8��Zi
:���yܐ�3��J����u���x�'�8�&;CT�P,�y���
/�wЖ�yG�YDW	�=���Q���G$��W���2�vT�DPqG����C�JX�$��#.җ=���
6�`�'9��}@�ܑK;���֓���>*�׊������ûb;����>�5 y�[�y�༭\C��O��&��;h@Ț�Ia�A��5Q��c  Db�J�״�0�_�<R�-��d���id}w8{�ՙᘻ�(ޢ��$�	�K�б��=��弅��y�?�Y��8�9����`������.Ŏb)�)
u��m�>ՈF��i�X7�c�c��˭�-�Vvd�S���4M��wȒg1�F�K�:�����셔��+O�f��}�����B:��j��M�+��S�{���{��o��ky�+'P#��[�����"����9�֍
,��f=��!�ROa���UG�����ci2c/��{H7��=�t;�*<)���OS��k�hp��5�W��"��1�Æ�BY�tc^y3��v�y�s���<���l��U��wΜ�p�>��\�+���3�)�k��AG����uwv����'�T�����O4���Ah��~��-xw��z�<!���q1�A��>�W���?����k�W)��v������b炰]��Tp!<!Y���:�}�Q�Pxl�~J�bR#b�-h�p^G͜t��К�y�P.�-�>��պ�o�����U�ˢ�ux0S����_�r:ÿNL ��g�bκ�#Qqsc��H�Y~�8��ㆧ�HO�����ŌB���,�&�3�DC�"�մ��� ȩ!J������t|{�0^�]����/bO\��Ps��tFj\�}�̭MoD3=��D��P�y�k����%���-��`m~��Y�cY�UFI��1G���tF�0	Zm�+�C�3�.;Y��v������)����lAp��֦_�ي�ǫ�Y��\�N[�l��_(pKp�X:�D!���[��fp�V�>B#��\s,��eBs�i��!�gDϨ7� �(���s4�ס����R/4O�O��*�MdK�S8�$G�h����RSI�"wr
en�1�?��뾪E�V�L1�ǈ}�x ��D��c`5�r�6|+'�040&֜QK�QrSd�nT�ᠵ$5ȹ��g_B�T��l�b�b�y��oe�t�C@Q�U�妪�!a��<`�
f���<3����ђ�T�h$0V���`��7y���\P�(!�c^���<�
k��VZQ�mm�5�M���ѮyC��a���;f������=y! �:�;4e	�'�ܿK�$�T��x�w��T(�������R#�C��D\�&4�
��#��_`Q�����7$0|�Ȃ`��y�Ntk���iO�d,
����a�_�*~��d��0�������u�}p��:�����z�E߭��-�D�5p5�sѧRԑ\�O ���/������f�"�=�ӡ�Fz}i�Q��wk
qj�����z��V��q��ᤡU�ɷ���of�7��o�i�.d�(��rĘ��1��1�ͤ��̞hjwTЮm�d<¯~k1�h�z��$k�nF&X}���;��l�(�S���ެ��U�\��p⽐��d���3��Z,�Hko`���2�W�$^3|�t�qx���EK�%^�;�����ژ3��<��U��Qa4ހ�^� %,l3_����E߰B�t[ WND3|�D�����:t����>��x=/4�<�=�٫�B2;78�������fcbP���bO1������//�L�CY��w�a�������>S��8H�����R8�|��77�gC"�48��7Ctܞ�v��ئ����,}��^��M����ш�����r���<+5?���M7�����@����l���7D$XT���Z6F �$��C-��)cK��/�!3�x*��:;���#��C�n�4�(��"������X%��ZY�E��p��3fŷd�ftG��Y>7�	�ق6 M*��vORkdI�%&+W�#����;մ�N�߭��e?��ߜ��yJ�%M#ѥ�q����Vc����Z��R�p��_����l}��^��H3jp�x�u5(LT=��^���i��ri]�!�2���5�RV�ŵ1�QM<N���� �s2��劋�!SV8`j�҂S-ISul9��Bt�\�����L�Z�u��/�J`���j��ш�e�a��)o~$��z�8,&�1�
	�ꎆ�Ľ�0nߡ9�ԤzIz�,�ӈKQIDЫZ
&��R|>����!��k���E E����2�(q�Q9�Q O_Jt'Qˤ9r��h\O�Aa����*T�lEn ]HUW��۳�M��F�uCQÄ�oO�z�8��W~�>,֥t������B�Nw�dR��9�l\Ng|w��M�9�������lG�/�?[�w�[�52�y���a�n�K��A��\�/��OJ���wX�WA�6֝��S�W~xX���l%Ր����]�s,����t��D�q:q=f��m����t\�Ng�dD2o�O=]�@�Go��4����KaE�T|�1S5To0���,�/I����J�G�Z�(�Į+i��7�R����+�1��J~T�9�~^'&j�2���!j-��/� GΖZ\��%�Hf���в|^b�y�{�n��j�'T�I���O�~,�P:g�+ǔ����}�Ak�������f����N4���1G���5o��1A���Jkٌ9m���+M�f4t�Tx������B��J[�}�����V�W���}`0���������S��K{O%���x�iJ���|'Ekڢ~�S���k��
��ݷ�(Ua�6��l�uY��$Hd��?�C�T����yq*�]����⮸�a��I���Y��OE�e���h@˾��i�ڼ��S��!h�_�C�ȑ'(귵?0V�����K���p��z䣘U�Q���R��`�����"�On�ˣ��x�v.~�h�Ąc�J����.^;��s�o��tC��|&S�7����8�A��X�Ԃ���6��^;ݪ�߱���`���}ZD�\?8UdjY��y�GZ��n٫L{��˕�q��D�u��Q"��\�(�&�1��Z��z��%�V�ѤAۈ��'V�J_М��~r�V�4�j����T��j��ˠr\�Yy>�Ά��%?�С�:��j��蝄�`*� '���S�Q_�*�H�qb�A��MR�/T�m�ՠ����R#���H;��"��Q���(:��8L{����}�d�T�f������9JV�m'�U�
�>�~���V�ϥ�lw�K����F�;(z�ܣQA��H�����l������^�� ��Q]Z
��~�fT���ޔz���ڤ=�`Vk�l���sG2����K�m�/�a���v����OI�p8hy�h�5X	���yޛrc5��(�qɻ��2c�e�
SV����<�+|z��N����W�C\c�����P��۹�'�����7��Wک��u,�����l�N꿫��읠!C.��=[�N5h�_t:%�;uzb:'[��JuI�3�VE�黿�Z �}-aK��@+ܞ���Oo�sɻ|���}Z;�5�T����À|�ә����|�1w�V�[	�x��c��>�EL�����j�۷_�N~���ȼ֚�q�{QWY�Z����[Ezϱ�'�0�_�C,aFeA���K;�����XZ�6�KȒR��kU��鱾�~n�6�n�,YI�qǸ� 3��̲��7*DM^?�e~��U�_�ڜ��4M��0hcV!�>��"�~�!o�u}�הĸE��G�s;���vf&&�ڹ�v���%�����%�gl,�4fK��c���(%*����c���
�B骧o�0�I��QP �s�
��6[��x�qmk�Ӗ�c�r�Ճ�Wf�]?��Ӑ(�����ȃ�8I�<:�x�|ɼ��9,!�L&���c�:u�3�ha_4}�2���G��PWW���I�� |C�Ϩ�ň��_^[�9n3�����g��ᵉ�ߧ+���w�'Di�3�����f�H)�V�0��� kM�y3��5W+�I�x��?�W�D:�v�������P�]��T#�k�[mg@>	g�$���甤d� �7'h���|r�2�*��o4�N��NU�;�_.O�4aaz|(��i⤐1����w�G��%S��G�9�T���G��w��m�����u��`���^���}��V��� SM>k6� B�Ɓ��xcJQR��&� .��+;�'�����00��׊W1e:O���"�C����<D�\���lM~���%;x�DKot�;�W�w[��*iL)����ƒ�f��.��hiX��4�{��΄��L̯xJ�Z2�^sIC�Ͱ�V�P����p�vwo�a��*���ǮZb.2 ����] ��϶�9d��x���`��P*���W��a`���n��9z�9Q%�H�Yۑ�^$���w��|\`ш'O����N��[ܯ��q�7�%�0yF\���_W߯M��F:��Sb�N�]�v��LC�iѡ|}e�,���_����f*��r��m�;7c�Z$}o������Mg����вk#f,ɔі�o���� �uM��YYm��M��n	.�~c�f���H�jb��WtT�@��K�H�^���*anY�ESJ�h�L��z�%�I����`ZN�w�@j,���֘^��-T�����V�WG���N��_�/�|hXT�z�-�ZK���S � xYz�F��ܯ�9�h�tj�������vU�(�5��{�Y�������w��X��1�㢓$�˵	A/~Z��?�&�_�zx�3��t Y�`�D؆LѮk�U��� ^�(b���Ck�����T��>�?{`m)�g4���3��4Pc�"����H}�bWM�3Zs���gx�5p�bCh���J��[��%���㑊?��Ɨ�ۣ�Dg����2��Fˬ�S����+�ne��:>��3rYhcrT"d����g��7���[���n���5D!`U�� OZ~=qŷB8]ք��S���m�&T�U�ؗ�| �Dy��l��[��ҫ���{ �ui�yA�KZ�����K*��Ŀ7�#��`q{w��x�r{�h����l~�PQ�l�;�J�\���*!��8�N�i�7�b�{��0���P��H˃��
�����O��k���LI2�ބ��&O�R=�?��BW���I���;X'�7�<��3�U�����Pɬ��kr{�+R�Q�"7Â�B�J�[��Lp���O�6 �}�Xs\Fp�uʧtS�`��dT�9<�h "�}T�ҳ�o4x���$�\��]��Ҕ�M'���d�ݏ96�'I�r'��{�T��)
7}�A�]�_� �	�t:����5k��P˕  nZ�U2����3%F��˴\ɻX�R�`L��.�~o2O�Z�T�}�D�b�Fh�ŝ����rw�m�Z��p�'���b��$������,E�.�?aC	���g䟧T�&]�Q�V�W�/��2&i2KZp)أtB���N���5p�2�rT�'u���;�K����6�7D�Uf h�K��wb� !��ˏ���� ͮ���r��l�$/�?��
;��oaXieEר��jr:l�)c����J����r�ћ͞h�L�Z��Z_?�.�;` �)�:�:���Ԧ��荶#��_=�Rmq$����g
;%�z��	t=ymX�<�rr� �u=s�[�U76��H5���.�U�����Uۄ�������M�r,����Tgn��`�BK��&x�pc86�1�.kl��:�it��2Q�#(�[`^Y�rd���uI@6���w��g<EDQ��7�1��%�B \�=�5���w-��V��,���|���S�z�{�NyE��u;�H\�W�����f{�{0�+
�.��E��P�'ф���F��)��[#�y��h�V9����p���c���%t��vtrz����0��0�;��� ���8�L4��@��j
4�hZ\KXn����]}>3�xX{����5g ? �e��H�!��*i���J^�������k��3Ol��3o���3���	/{x��VY����G��5LPe)�h.�^ �lz�sx^Y:5D�oi�T A�	±�	�����rt�$8C[��D��r 2��#M���^��(���r>_�
BQ�� �nll@���mm#*++���V���&�������<!��2��d�i����&��z`�Hl�c�y�AT|~b3qC�.d�WT�`����8��~ �9abI1i��i�6t��ݪ��;[��S!rXq���w5}� o�!���#ɍ+��@OO�6�7@"~� ]����D$m�;�R��N�qwEG����6RQA�M5�l	�Bc��hf��L�����h�q���$����b�Jt�R�O��l�G��_��3�+fR�����(E��XJ�1�Y#��7D����"��g�K���tCa}�����OÕd��A��/��2)�	z=YX*�&��t�F1]�a�6�dٍ�@|V���nwÉ.�Ԡ'N�`?�~�.K��[J��P�KM�k�_!����K��@vѵ�_�@b����_j1����xp�
��p��gSZ{�=�'~�$��Ƴت2�B-���xZ�C�
�0�ȝ���ہ�%ηe6Z�-B�Y�O�>�R�gg݅���܊��+�E!Á��e�2���W���1\��xWgdW�K/��H�_Q�^LGs�� �G<%��/�j�ب$d���]i�/�FS�My��%�3���^%��Q v�!X}g�<�v�������f؜�D�7^)	�K��1M���ZC��jC��iC-�h˽�[�y�� r�ߞ�/(�+ף����öa� �2�j&zL�2$��~�7w��J��V���
_6��Y��,<��`��)���G���f_�,��J������h�<����B0>Q:�S�$��
�Alz[|�>.p1E����� ����q��	Ks��TD3�b�����Gt=��`����b�Z�y�(���qY�R�B-0�h��9��0Ci+?a�^_�Q[�[���p?F��qj �s�I�g��i�٫ۋ���C���;`G���8�j�:�/��I�b��q���ҋ��@��5ňZ=M�T�4�-`���F��<I���D�%�y!Pn��n�7���㩩�ubG)�t���зYQY��(l�E��M�C���(X~2��bY��]����s�|�A&6��V�~p"�!z@�!^����튙��j�;5��Q��_Ƅ��6�����X���"�����S�pAL�9>q�����;��`��q^�QV�<�� �6���3Lb@��<w�c��aɡ�(�
F�� ��~��?Q���`}k����m<�0?�I(FQ҇W{�ꥉ�Y,:̽ CY�7��S><'��waI`��u>�0�©ݔp`��m�Vr��7i�]����J��J {���:�M|��g��pw |�VOA`��^YU�?���Д;h��AJ�s>.Θ�� �{��-���x��t�g�J,>Yh)��v4�?�Β(��-<W�%���T�@ ��c��+N2�qPx��*�N����B��C�T�+�D>@'8,3QW1Є'p/-��#}H/$��;*gG?vFm�|��/�����񄇇G��I�q�9(F[{{��Ƈ�fz�?�"� {���Μ�����$���xé�������h��ϛ2��J<qh�[���ɬ+n���׊@�����7�M�W�S��e��A�Vf�%A�O����v�[��������$��TʉzN�"�agyx߿S����ZOλEr�w��+3�?e�H�5ҟ�9�8�O.*ܦ�v1.���
|wp]�֯����4�������Fm1
P���!Eƙu�s����Ҥ1CYT�;C֔ ZK՟ˁ3��.�Qۊ~&5�B���_��a!���\����a/��H8&5���3a-�,�̓�U[w� !-�Ggw��L��cv��'�ѥ���������-,u�m���c3�t�&ْ�l��r4Vt���o�B56_R���<�"{���4���D\i�K�~��!,È
���s}��2H��t� ��+R���_6����N�q��W�!$P�@��H�
pT��V�Ds�TC��'J	���.R]7,�p$��h���bâ��J�W�T�Mgg�<Q}.y��"�]m��[���>ͣ�nR��,v��]���\�-�)�Q{)�Ry\�L�v�#��W��T��@P��
��ih;���.I��؋�(K�U�5M�S0���ӓ�ѧ����'��n������Tѕ�c�R���o-�|h})l��mm|�G?���444x[E1C�����E���� I�X]�c��F`T�����5�3[Om�}��*�Mj�홠o?i���K�Κ�̏J)A��#o���r�ߟ��;�S�H^Cm��чM���6�7�.��d6���%�ū��R�G_M?��L��,��U�,�ކ4���v�.�a��MAl|C���VK%W&��8NB�/:��w]n��������z�3�4�����.�b�@Ոj3g-YUhK�TVt
�����W�no��L�d~1q� F��~6>{O��V��Nw���Q]g��"��"j�H�J ja����j����K�-OàF���=覆����I8T�H.��Gq�N[H䧓	�*�aG��Lzz����i�"	�{T�O������tP\"��y��W��Q*����g�J�f�d6G���P
�U�ʨĲu�F��N	�Ƞ��LB�x���Sb*^�e�I�)'�G.���6�����Z/�*���OW�,�������+�Lma�)��q{���[vt�5\U�bY��b�����Z���.J3H^c�c����t�zr��If=!I��������g�%i;�������/��hna��K:�듩���t�����~�_�gNΔ�F��w����i����B�߼׆�t�w}�(�3����H]�@���y�P-'`�<�2enxAU����Ϩ$���Q'	v�ihǬb��ӷ�����6;~T����>�����Y���ͯiP�CL� U77����_2(�&��c���>�pFz������/IĸY���d��p�/�(�]1'bZ��lZ�M��YlEj��3�^	�G�}�~~�w����W�?ZB�}�V�G�BoȒ�sAWL,�+q���f�����ӄ*���2|h>� ���Ѱ'���gh'.��"Z�z.Y�:��q�A2P �=$�u@bi0;DFv�"�~���'���|ׄ��C(��]��N��?w���&��0��:xpO�{7�Úb��4p��`�ɤ7=�.��l�\g?G��pBg[<_��b!��Y��옽1,��C��g��tv��}��~�����qq�p;����!*���z�vC�(��W#�)_�IS���9�ly���Mi��W�[�����x*~pu�0���è���"��DDH�P�X��N��D$|�'������(n�������?�����7����fI$,�{4{]TzD���e��{�4��)�����M�%k�?N&t��6-M˧pͫf��ܻ�I��.��5�9>EB�}���N���9,zN`�� ����<��������.�\�KCڗ���m�����H@�z���|��ĒfǱU��n.`�0�S�Z��;����y�>�F-�'�pɻk�E�;��m��n�A7Z������P3K��0�ػԑ9�w0����������X�҈�T�l���l�z���>�)/�w�d 6�D�ql������&�cG�'a�B]�mJ�����8.)Dm�P�:�|ɔ����r���G}�\�@*�j�1���,�թ��$�1ნ/�?�79eJ�ƯE�������v�`�$��/+
��S�֯���9�4�5�4���aT��,��}��=��	!!�Q
	�4Fm�m�H��3 �C֖$xs��)oj�显���:k2���+!j��T*B�
6��-�X�k��<
O'f�Y��K�Fޝ�4�t�e|qo�gG��b	6^��XU�Y^�׽�lo��F��EQ��P2�����l#;d���(�6�b�5��e��eo(Gq5�Uv���w}Ol8�g
C��ep^��霑06�@%Gu��߽b �F��h���3�x�4z����a��f�$�����U�sd�Ι"�pG1Ĵ���K�����jd�UU=[=p
����6c%����;�(��o��m��[v�ף���[v�W�.�: a�k�E��?m8@��W-�(��F6C��ݧ����m�R)ά��T�N(�+	���
��������[e>��Clߗ��������A<[h��c�$���`ɵÖ�F ������g�%��U�¿؝:�:��Px�߁���p:��}��L�����#����� 0X�����ܥ�eߣ�`�Y��:G5�p@��3�1y/���YB�:��׸f�S˾ȕ5-L,��}>���Q�,�B�;ѿ����6V�#�a ��"~��w��p��Diu����b~[3��m����G�`^7����Ac���,���s��\���}L���s���|mfR]v��4�>�m�����7?y�<8g��Fy�K)v
6Xc�B�d�R���'�Pi�q{p�'������|Iisw˄蘝�M7�ŷQ~0����Y;�}n��Xqw��
�Q�0��r�8�o9�5�á���F�<��>3D���
�-Ka-<0�!G��oC�����0�Ƥ��(ٹ;�Xdo��VWE��ZQȔ����[��&5���md���J~	��귒�����	G�@ˇd�f�S�I����1(�V�tȁ%�.��T�"(Q�;��#��,��s��n�lum�f��E�	��a2X��1I_4Ӛ�9xъ�>xvR��"�-����.��QW�{�U����V1��F�]�������H@fTƬ�U3�aV��#z=���b��tS��ۈ\�3e���+7D��9{ߺ�Q��|���0�^�u��af����v~`�8��Ias�W����aYʾ�v��H�Q��m��&h�ɖ���^У3K�p�fr�����v����{���.��v�0�Vd���,�(�q�Ϩ�ģ��P���_�Sև2Y�7���#�S�=M\Gyͨ�j�L�)ڜ�q�-�c�5~��x�A��&�s&�?
�cGSvFu�t�|mJ�mAC�}ڹf~�͊`ry0�hm6�>]��*V0z�A���򕗵��'��`��V	�6p`��=J>�n�3�G`���w��K�2O 5�]Y���hr�	�h�豱��`���\G���5�,⫼�DC�IP�]K����T�}��U{�pU8Ma�Jv6 OdH��
"c���[��� ZO��|LZ�������%y�+�l�˃PK��	f�ןl`�B�S�����{�Ⲍ� ���H!�m�y��,���1w��3t}/����m�(�@�03������g�R���@˨�&%�4�zi�C~-ib�ɡ�û�A�Ҟs��O�V��q��?�Qb�����5E#��1��)L��%@�%7M6�h]o��&�Ϟ�q/�ģ1���_+W�h@�cW���	:��!���}9���F
�̶Y~*�OoTT���8{���"=�bI�H���*B���AO��T._�g�Z~�^�)�̣�0j���b�.�=P������I��� ��&��\�%����Ptώ�Aw����ĿK� �O�d+)c��uyT����7�4�<\_E�[����M��������J���b:��!P��h�g�%�[6�e6@9�����*R�7��=�yR ��忊�lx���/{ ����i$G7!6����SD+��o�:Q�����d��
�h�fW�W���5Y�<�k����W�S��m	�V�$�r}�-c�j -F,t��:�kp��U��6#vpf׎k��M
4�^NGГ&,���/�t�-�.�)a�=oy/N(^CP��X�Jtޥ�w��=�'��`�-��:����8.+٨iUt0m�8���v9K.����k�e�2V��{�/�Y��I[�%/���t��Q8"2jh�FI_V�4�(z���#�~�OR����=]���r|$J	qL�p��usu}���~c3D��o��]�2L��������d�RRz^W�j\��i=�+�t�8�+�L�m��N����FY!I�s�A�,�rp��f].�]���9OWy����� ���s���o<��/>ίe|<��>�zy��(�;�%�X���-���A�H�$63XT���$�_�19&�@ٞn*�!��dep.�vݽxpMg�o^[���^d��i���=�g_��WVG5�pDX������?Y��Ud�����-���Ű����lf:*�XA�"�7�!kZVQoIm�B�'R��)�^C�\��'��7��"#��A�*�O!�ߎ�i�o=5�Զ{�#�j9Y���.��K��O��m��#~HX�mWTJ!z�IFľM�V�My�@��v)^�_�� \��̃���kqId+
�e3f
�E�m4�ރ��������4k�L�懃Q={j�.��z ��+��$��dw�8�^ڤ���e�I�f�q&K�~Wh.K,��G깾_ka[	�����g+���0��l�^�τ�B�M��u���tL����8��d���[Ӕ,�?vXM�D�1I�k�:�&��
S�(�t����m<�IW����h�V���J��x�D�,�L%N�Zr?_�`2ب,#k�cqw�݄����k�z�d����z�LQo8�qe��Pr��3���j"]v����"D�"�Af���$���'�$<s�3����/e��kO(1�G)��Q8�UK_�I�5�u}K���)���=���.a��K�c�B�6(�/��i("���r�������	����'=,޿,|�vC���1��LJ�4s02�7Y�!Dei^���3��l�s�A���i*�t�nJ�^����l�+H��bp�����H_�뻆�ؒﱸly,o�VEn�k"|p	</�e����?)O*�z�
�s�kLJ3��׷w/�<`���b��9�C���7�g�_�"��H&�}��ݜk�����:ִ�_�~3�jf3Bye��	�#���{�]Y|E?Kd^�Z>�Ȼy #���[X�ۡ{Qסr���m\�TIS����f��N�ߏ�B�t~����09�^K<�8E���I37�s!�x3?� 㱿5���$D(�UĒD)#��@Y���/�����GiNc�H�ȯ�TcRB�r�#yIoO<�h4) @'�g�~����W��r[v��G����?�pܔd���똆�Yt�6��/;�<U�����!@�/�[�����u��a'�����;��ު0��b1Ӿ!�d1G�xe0I�������d���1��H���x�[��Ҳ��+l��CJ����7?�;��[/1�R�k�^�ڈ���������޿DDD$����.��A��Q�nTr膁�`�������x��w��~����\s��s�u݋}���zO�ך�}I˝�ׄq{�&@\kT_?U��Ai\ی&T)m
������Ү��p�7O1���+�g���
��G��0^��r��@��eY��E�����H�;�(��J��Wq�Un(�l ,���%;U��ַd��Ш�$�5�Ml��#���I@�i�'�]�@�0��%��ft�8������^z<�W��.��z!�-T2���#�
��P���ڒ.�%o}u�s�\�Y3[�F����1����#�Z�yM�އ��υ���CLVg��FS?k����b�F��޹)���J�[�gfFt��r����8��L_&�~su`<z��3��{H�F�-;�J0~"��{��q�d�V��'� ���=��o|U�"��	���ea�ɭO9�?���J1�fjXhC��'�/���Y�;�g��
q�.\�m����w /���Ԣg�`}��ad�&ߝt�2&��ۆN�^~��ղ�k��MO��\���@�r���8*��l��V�y�����c�c�B�F6/l��~G�à�h����X�qta����4Ve���K�C��Y�;�y���2�5�@[�Z7��=U_���˶��%	���������A�J�!C��Cg-���y��G�P��E!Jm���3��a�3I��|BI��Z�&$�Y�o�x
�T���Õ��������Z��G�)�
�j�r�4o��5�t�_���~Z+#���v�I�y��S�r{Y��7"J�bU����&�Yc��)F�j��񇧞=9��+�W�=�p�iЬ�fY>�"s��>3QL~�7�� ����g�J�>@��W��m�8�TT�`��j��Ҳ�lOƻ�v�������/�qv�=Q��U��Sc���ό�I�}�k�w�t_�0���� 2�Q��W�h�k�=��n�0B�)Aa��B$�� Z�l������D�j�3#xi�q��V+��LU�Ic:�a��}���v��/7��Z�s�~�W��)�����ٷ(a��O���r���72uO˵��y��\ބ��Cf��������H�)K�᳑��h����F�aZł������k�iZPI(�,��=�՟��* l��wD^��݉	��Đ��o��_���ӯ2���^ӿS���{W��w�\�`�����dG��˸��BVF��O�AJ�9ŇݍX��= cz�1��&O�s0"������)-I'�悇S��~y�XP���39���ptk\4&�Y�@�'\�}�u�c7�巳b���"u��`�,z�'���Z�(�]�;̀�hܞ�8"F�����]>�#M�ȌhtН�+��i��w4���������]E��r�t��a��^nel�m{��o��VE5>�f]����?��Oh^��f�}�=��d�e�������ٴ��{�"�eS�¸#=�l�ϯqK$�j���� ����'�~B�5w�^��@�"��>~���t��DkM�Z*��e�9��B�SB�Nl(����8xb��<�{+����y��w=��:���8�I`1��բ`o�����$ȏr�$Ii�1�k���7-��(X}�"QH�Y�f�U�m��oFH���ӧ���m	2x��y�UQ)�<Yw"r����9*��6Koj�8.�Y;��A%���#�@�a���"��,H���ËըJ ��I9|�lqq� R7�O�+�ԍ{JO���c�K�2�]�uqЮ���3�:����7i4oW6=��%�9��+yk����I����������";M<�qV���dC�J֯c}���F�~�J�D�WF3\c�\O�rÙM� �b�
���p%?��u>^݊ݘ+���;����r/�2�Gw6�"n�Ef��=&���)���M~cάۮ���e����l˺��C�vm�/��\F��OVk�}�
�����'��j�M�}k $u�8�����9(���T��
��`�'q�*����B�'�Y�jNe��]Y�ʶ�	O�'O��'I� "ZUV��"�dLb�*��B�х��������q�ߊ�sD��jrS���	L1(=i�Ia��5�/�J�ړyt̰�Oթ!��~=��������s)���[�w'��gU��M�ߕh[���ieՑ�Z��2�r�y���b[g���� ���>=���k����Σ!���ϱ(~񟴽��,�c/��b�ʯf7Eh�.I��6�������[kJ
I�C\�o�����+�}����?�_`M��GO�|�K����/���"ߢ$�E�Z����� ��Ug`L7�~�
���~��o�.��9�J�\�	��z�,bp`E�^ܚ�̵b��P���P��T�cPe#۱����\��^n��g�W�Z��X���?8B��P�{��$6<�SoH�Q"���Ƶ�7E'�g�jl<I+l>?�p��U�e�0l��.���e_���gH=�J�y���w'�����$���T������d?�ůj1G�)��8�ds���f��gtJD��Hk\ɽ&�»ֺ�� ����h.J�B߬;�;����\#�U T^Ԥ0���>#dN��2/:\w�����p��׃u=�fk't-��I����/L2m��]t��:�V�(�*��p��K����cb�'�J/���B-�O(9����1u3RАJr�I�2��cIKx�KZ-�~��B�j�tt��?Y��v$q��	��̎1�t��M�� �F��ە�eR�aNho�E�ֶ���᫗P�1j��'��f���ȅ�?�����4+ݘ�~O
�
��~3/X�N���,juc�uj|e8�5�?k"]>�ͧ��x�N��3��)�q�]�]�37p��(9_�Z�om׻F�b��v����(�Y�Y��錳~y�Q>����@E�]v����6I7w���{�L�RQ1�=�9�.MAn�-�X�����~��<��`�)D���j��J�RU��p����A���G ���p��{�A�X���C%��P�a����.���\@�ҸأIJ��j8Di+Ms���]���*#�Z���S���fmptz"hp��m����y�QN���m$E�����՞�7g2l��}�#����Ak2�����z�����ߟ*�-Q��@~c�X���z�@��i7�֛f�����yڤ{��d�?W�$1v<��sp��X���=ۏ�y��;�g)Ϋ�m��(+/��L����E��](dd�a���?�U��D>�Uc��n`}�`�2���߬7��cu8�g��i��悷�JX/�U�P��(�������s���߭��N��YX�����-_�h:��S�j<Y��o��[�m7=cL�"��	ȍ /F����#}�a�򵱺��fI̎�6]0a?l��ˍ߯��A��������3.�~�lL�/U�^�k�kP.�����cx���/0fh'��	�=yt�\YM���Ia�$v{ ��e�i�|���:�<�I�!�`�E��dV��Y��nk��N��J�f��H�`Wמ���ĠZ����mZRg��QLE��hlfqi���QDz��V#������Aox���T嗎��}��t�%Ģ��r�n�vp�G4L%�>����DQG�oW���F�����m��i�.��E��E2r
���@�Ֆ4m-Rx���<�m�
�ݫ��6E��^�/_��~�#N9��dް��N�rjn�͈2�2�b�ڸq&�w���.��оoج�4�Mb�T�3}�"�ɂ���HrL�W���n��������̧�.�|^�x6�wO[2�J�^�|�sx��r�.I<.����	�N�P�AGŌ�+��wI��J`��VjF&c�E��s���{�^�~a�_�I?8> c��8m�\
&~Ⱥ�.aT�m�sWG����Fm���DH��;Uv� �\�7���tr��R�,f��mr�,�^ =��l�w�^���nD:DCGI�AƧ?�� �B��S*ݥ��U'�,�@*�^$��LfM�Մ�ǜq"�n�� Sߎ�_)t��>S`�y�8W�2�H�����A���7M4�˱8_�qB��ƮT2a�(�h�*�M��,����ȄEY�3B滃��TAf�d2ws3)���I��d�TSgV��Ys����)]U��D�@�7>����D��VùC�m'���1��(�ƥW3�a�i�G����r3�D^�G�Hb����E�v&ߨ�K�$Q~۲-'H����(�z��U�����=b����ѷ|�+��/���}#q!���#װ|#�P�r*�y̠�>Zd����v�g9��ػj��-H1c;�;l��v����ތ�C�Z�:�V�w���l(��=�f?+R���O�y�ٞ���S3����2�W����|�b�Y���˽I,�|Q��V���wS�v*�L�ඪdr�
5	�{����t�|h#�:���iʅ�����ݙ��4:��|I:n���6��&�W}�r�@�l�D�b����%(�$6�fs��|��k��b��4�D����~Sg�xm,�q1"U�W>��Qz'�,��u�!U�B�|���{e]N��p�SCwC\+������f���Ʊc���Q��;X9�ճL��aGRi�IޞLs&���P�emNd/��([�^���r�'�n�&aQ�%�W9Q����y�j��Ę'��(&�>�3Kg	<����* �����ИүW����GlƉ��p	��de(Z� ehr�������z�����QbXx�������+3#�[�q�]���u�8��L�$f�B�"��kE��(D/��>�zM�PUI~:�\C��R#�A�����V�C'6�+�x�+���ÒI����Y[���8��;�k[3:��J�����N�?������W��n�'����#20Ay�{��I�/�s�3���K����e7��yF�|�*;e�7���
h�L}��D�k��^7m�V\�� �)0.$k�mB9K�xV�{����1��%��U�N�A��
pϷ��SI:qqե�%i�S:�_�!��;Kt#�S�M\�<̣r|bZ"�(��W�շw]�7ʰK%���7S\B�jX�z��b�"	�;����}+�UV~7���o���g�]���p��{W�^[ۤWz�J,���r8�4̙��)\T�zA��H��>�r���m���������UG���w��\�ס2`��)4X�ϴ�tY�(����d9c��<�8٢,�Gq/ik92���zI�,u����ډ� }���L�G��=��Lei��*��xW�N��+��ݢ/��A=aN���R��o�?�G���Y�����'��'b̺��S����,�j�O��s�uX�wG��?�%���F�s����e)�e����`hD�����L^�a��D��?-����x(����!�ب�w#ef��P6#�Y� ���d��:u�Ƥx��5YL�*p>�G��ջ�ȧ�q��6u�SS��m�gnDM;�͘O�!@��*qP����F� ����ĝ��+�2c�B1�*vo��v�L+l�Z�e*I�RgF���!DhY���O�4L��I���2R�X�fZφgx�(��Va;K����o����}�D��Ν%�J~�/ ��Ы�����J��	�y5���:���K�/((@<���M�, j�?��6;�O��_s��9�M���fN���1#%~��Ϙb�A�,�:�^�a������K��{| }�@ sra���5�̺&�����}q��m�+}����r��~���W{}�*�ӿ�ҪGG��J�E$�L�R�'��"]��Nee�[|}�Z�gOE�J�3�$|����CZ�L�"�ܤ��d Mn360����
�@���4n��rQ��ɣ`}�)�ׇ�G�震}Ua�����.Sa�l��V��6{��ǻ<���Tjg���Z�_::z������9�L�{���Cw�m�����7A��#�`$|�
� �����w���,��o���@z�7]|%m�n�[��ⅿ�L�un��=�
K�q����s�!�������8��?7�Q���)í?B��|�_a�t>�����\���9�)���0��ۙS7Ƣ��A���i�59����iW�;|�>bs~��7u�L��Sr�$W9�����o[�C��a1�E�_S�z�'��U���`�%�gqϗ �������Uڛօli��|V��[2n��E\�Ьf�8d�؃���dQ�JG!b�c��0H�y��=��z%B�|��Nj'D�����V�ܖq^�NqypDl������(Ty����y��$���z�������$���C#�G��*�H�K=�/Ka���L�r)�p&��e|�<��o{����o^>���٦��Dl� 9��K��V���v٤������l�r/��0��5�D��w�(�L�O0�4�C�8��*��֎1�����jS0:*�x�>�na N��+UK6�}��1i~����RhgqJ���*1z���}����Hv��J�)�أФ
�1��"ʈ6h���ͦ�)���u�?�_�YdXJ����|K-�]|-,��o�'DZctSg�X=��g�x�J,۳&�	�WH�P<��Jp߮�/�	)%��8Ќ��~Ȏ�(��ٿ{�� �I��z{�b��N���J��@$ҡ8�SyxV��CjK��U"�nF�4������
S����eA�R����L��y:�m�ٙ��E`�.�b.v$JxF>w��eÖ��y��R~�wN�����Q��Ma���}�R/G���Ƽ� 9�ك��������F�80���r���K�+�B�>��V��A��m���eL��3B1�d�Qf?��!_��Կf���f��9�����9�N I�����\& S�8ɻ%�ku��1Y�"�d�`��7*D<�Nsߢ�;"���S`�f$J��&��)�v��*^*Zz�E,��Qڋ�d���5��
oy��l��V����Ӿ��@���U9\�Pe����-9��縮ue�XalK��]�w�O�zd�O<�U?�����h\GMj������8Ѧ@��SD���&\z�����F���.$�I5L�Ex���u���owb,�kn�q�U�@�(W�8}o�*��_�Mz������'R/ 6D�q�p�q�n�2�XiO:�g�U��f�e�r��/�zG(ǿ�Kʴ�.Dtu���tT<�l���8ve5�q	�@�#N�:�nq�爗�ߜk�O��0X_g�lݩ?�[:i��wѱ5�,+���P�����3Q��0���Lg� i�*d�A��\L��5x�� D���Kc�2to�c�o��`�� ��iD~��N��:�Ϋ����bT�O�d���;z�Y�v����Vj�x�W���&m�����Yͱ�G���� ݍ	�0��!�Ѭp%u�����`8x��夨��f�lUX>�sL�<%֎=�fQW2)�H`��P���z��ܲ߁�(U�)����?�z�`�F�`)��ul4@�ّ��B;�sx#���a��)��y��*�ts�I��2�t�(��,o"�Z�����,�t��3
����+;��AS��Y�s�9A���1NY��~4�m�eK]���Hw����G��n��d9�����~�_M�^�U*�]&a���Y���%�u�0�Ȉ���F7ݩ�e�qP���xߥ���Z�>����O������JT�V��,6������d����@�t�F�{ڲK��Qi/��Qǡ��<]�z�ق��.e�9��hJ���w_A5����(:~1}��{�m��Lw�o¾���E���[4xgerb�ǑѼ_>�ي2��5Q�/�2}Xƭ��1Ypز�]*��E�G���D�Mn�7R��)T�_�ê��=(�����˄��>�Lm2o�]�q�)BX����p��n~���N�n�n�O���1�qP�W�7S 
a�7��?�#��B]<���sw�q���G{�[����3y�#8����Vt<�R?�XC�=yl�m����֘���L����|������]4;���+���<�C��\e�p�NԹ�J'�o��>�k����ş,�{dt"1���ٽf@g������0��"��6kA<y�U/dg9<!�ٙ#`��a�ې��������2V a�9dG<��,e�� ̩�Q�|eԆ<�����)�"��h�����K��9��ȾQm}�j�b�Q�����'�ǯ���;���d�>�3�`����].ي|��K��oݘÕr�Sܿ�S\X �O��,�e���zRo��4;$�ר�(,����NL|/d�y!z�9X�H�ш�j��ss5���i�(M&ٟH�������B�z�%�wM�zl�}BqZ����J�8�[R�u��V{\��V�|��+��9A���I1]������Y�У�1����� ��K���ph�����$���4�p�m9V-���vخ���٢`�!�3u�����$�|���B�2SI�Ӵׄ�"���\�����5�ȉ*��.8R�֌��ӗ?��"�L�b���96w�C3'�̡q=Vc9T�ڤ���_e��s���剷B|X�򽺯d��By/���E �8k7{ z�qt캑�1�w�y��f+�Q;����ࠑG��!�������`�L�Ȗ�,2��+�h`���Q,�� �J��!{��@���C����C��D.��I=1���սCcl�gq*s���j�H�.[�`������)Zu�"g��k���]SJ���*t����5�ֽh,�;*D��}��{Nhs4u��;����q�'�p0����꩕�c���c�abi4��CB|>`m�����V@տAx���h�fhA(�B����k�g�@uH��d�4��ϛQ\u&X�:�\��AF�u;�)_gnXi��:v��$�(!?:8�����iH�G���^���u�i���[Bp��w&��#��!齁��"�o�%Upg��R�����mT`J����aP�Q1�C_d�ߖ���F�)ht�V�y�I:����^Ķ�xT��m������/ƺ�gv��c�E������]�!N+�li��c/��2z��vq��I;�R�Oa{L����5d��ơ8:��U�l�a�5J��E;�����.�a�X/[�*��h���CX�%&��
Q�Y��<e�tm�P��d��m�z�{m���j	�Y7��Q���Es��m��I�Y�z6�f���M�V��z��<4�^�`t��y45s��$-�W揑Ÿ�����9��{�M[���a�/��<^/LY
��[eА��sR5S1:˛�O�n���4�V��
N��k��g�G�"{d��>췏��$���z݃0j+�d�2�*�)��d��Vu����nu�3��I���u|!ؾ�C,G����4c���^��Wn��p�+��Ks�YXג��pѓ^p��j�`c�ki@�V�#���{�f"��fL��@M��U���"��O5a�&�[pH~�N�r�Ds���]��+<�,\2qy���u��캦�ݫ�*����Da�eI�	r��ޟ@�@����E9r��,��C�k���
8��Ga($��sFZm��9��%w��`�� ٣�-j�=����4{��G�	�=�2�m��t���m~k��=��Y���T���`'�w�4۬��n/V�sg:�Ǔ������cn��6?�W$Yv�0�{������^݂�ݥ�{�vU:�\>w:_lr��G ϰ6����gν�}�j�«�7Z+�l�3��]��c,�&MD"E�u����10zq�7�oJL@;�},�����!F�M؊�~����� ��O�$���F�5��P��*Ŧ��B�a1	�ry]v}��[�j�I�t�Q8�/��-9��f�$��d��Ϝ���GAhOO�԰����#�dh��nI�o.��q�VѲB��׎����>�N�U��:_Wv�Љ��#)G�2c|t���_�V�2���Հ����
��ݯ�:xrwB~W�+�>��IOT�괉��@��E�Z/���FT]Rݤ@}�i�x�H%}�Kv�i����FT�\-�s} C���=�ߜ?NV'Lqt�RE��+�@�/��������QG
������ԣ�`k�����?*y��	!m�wݭX����)��-�G�M�J�3���N�q��	�@�B����mµȋ[��,SD=���}��o[���z��XY��6�'�������y���� ���������K"`-�T�ʹ�\�kﬥ�m8��2,(!,z ��\M��n�������(���A��@c��������sWޟ��X��VӋ��#M6��w�V����c�!o�Յ@Cא��/�nB'������t�i���bg�m�C���ZWgq}�D�Wm�]l��ThI�X)��o�m��;&�vt9v��!��ށg���4��>y[�9�È�w���]�����G_�%����J�Z�2Go+)s��ߒGAHƻ�<�g�����Ǡ��2X\6��s�W`c�S���w��oZ��9��ݿupA	Q������3�5�5I� ���^;ZY%��z:��~5��L؃���W�~������^�I���H�J���j�.�t����D+�>��Wf��'a�9�� �7�|��qշ��n���Y���Zrg>��?�<o�*���-�c�@��}'�;�ˌ��F�70�Z��
�c\L�)h����)�`�ձBwk�Q9�#uSU�<5�WOrL�M��������6R8; �UBO�,�ܛ񃬽u���5s�sa���������o�,��)��/1[�7��I�Wϱ�k�Ʊ8�7{c5fI�=�H!fYi�u�<�Y��R�I��[-�T���2&���a��c�1k��w.�u@����m�)z�!}�>gI�%*TiS��pZ�x'���-���S:b�,��<6REB`��XP����.6%P+�򶈗y���zTv1��X�Uq��{C(Ԡ_����g�� #�vf�åL��<$ί�T��ͱ4 �5���q�g�Xo� �x?�d *汉;#�e��T������z�=Ke�Dp��Tқ�������a��\� h�TKg�bS��U�	_�W�N�
�G+�H�>O
k�e����������_}���4C���
��L[{D@N��U����U��]���Ҁ�� 0Mdy���7���ޟ�-�}7�/�)�qzV����(A�.����ۂ�m���`6/�V)ﯿ�f��?K:�� ���F�_�|��<>z�X��Sr:~�?s�������Q�癫��3��9�?�@)�bWU�;����Bu��~���x�����֮\��ָ}�L� o�OlKp<����)�@P�`'
�&�ïBr�Af7�[;�2X���|\f�ľ�lycS(F��o�O��q���4����2m��ڑ�2���%�� ���5eL�^谢�\�q�e�Q�8�Gv�����D���pѤm̈́�}�[އb�9Ȗ����%\eOZ)g�_�V-=]�C�sr*�q**�5�(~�ٜY�AW��Z*�;L�8�0;E�=�^��=�:�d ��,��W\�J8s.Nm��b���RH\@��`0���z����x/滖J��I��}�J�`��I$߭���[��4����A����1�B^��|_�գ M��}[��5���N��c��)�y�q��%���_p�j)�+L���GɱUtͮ��ou%j���Nw�'��DM�,�}	�%������s�Bڒ�?���k��`+XiBB��1\'RKz۰˔*��0Z%ܼ�D��n�TIG��~[��x�:vm�04mM|=bK�F�u��{�a�~<���,�Q�gV���P��{�V
c�53Pg���ӳ�F!�\�
�C���	�D��N�}q5�eO�6�^��n�Ɨ���%�ߔO���fn���R���������c~ Eܤ��i�j�k���m��,M�\.���g��(�V�r?��	�3����[���q����ى�!�6h���@��,;LZ��\y-4םn��	Ux��:��C5�2�4V70O���3��x�~�Cj�~
�����L{
2P^L�?z[�qO�Ƕ�gso�UA��������p�q8��h�w.R�����}�\Ƥ@nj~�G[��S^^��~��kX�~9Ϲ�C��=�`�ܽ+�Q T)���Sƣ�L�gud�N�3����p��1�(���0${��$��Q�0wL�w���3��Pg�X16
����Qlrul�����&���qt��k�(J��2t�s&{"��,
�?/�bt>b`��-6 ��L�T��pK���v�x�w��ƫ�^{n^w�_�ɼ������jWU��PJ2�_���x��p	Hg@ �\���*ފewD��wA.�Y����������1b��Y���r�mؠ�Q!�w���9!y�WR�]]�4���l5�k���.&��O3J��������zs��m�([�s¨��N]��]����b]wu�����.�A�����4m�h����Y�f9�>�]f����Y}��dR��ݜ�;�Ѭn읙>˙ܙ��5(�/�G���s.E��}�O�����`�쏞l7�u���=�m9M׿�;��g~3P���|:N��[`�Uy�` ��<�5F���˗�D���S:�������(R��38���&����:�(X�c�״�r���b�㨞��p��q���r�i�]�]W�6m��N.fg�_����e��wKCQ`��5+��I���Ӳ�_�4��F5S�� ;��|k�L�kɠ�$N����g+�_[Yw_���c����P��j���M�kx�a�.��?�&�4eg}�?�%�!/W@��;~7묞��.�{H���xgG=�����H�5�t��f����gIh<_ťH�p
�,��ǉ�l�ߺ�ZQ�W�W+��f�AP
$�GU4���������1LW����]@z�\�����Fc�Yо��m]�I�b�<B�ݣ�`C{��l�talc/W�k��r����ڣa�ȯ_��.�VA�o|�T�R��]+���^^���R.7����NGAF����0p����~O�**�p�6KP��bcZ��ľc�ݫ������&}�>��5%�&�NG�A��"/�o?�zSk�Y��,^��w	H�O2�pF���M�B\>�9�t�<��X����d���Q����6ܾ;� �I���{�;�s9�t�5�X13(I�򎳶3�W��I,���}$�Q-V�������n@0�~K=V�o�9��N��p���pO�����~Uie��έB�Ϫ�n��[5j4���
{�$�<���{/ ��}5�
�1�����}����ߘhFR���~���� "���]f���Oyzh��܁�����dA:f�&�8-�l��U�5+GW�Ŧn�ǔ�6c;�[z8���У��� V>$�,�!,ř$���p�H{,ǭ�
��Jߥ;�QקV:�ȮԎ$�G}��#Źy�MOgm/j� �fe���~��ڷu/\�QYI�f�0<ϗlҡ1pԧc.�\dCEe��`"�_�ٝ�?�ljm��U|l&�`�������_�O�
w)~�!K!>������{� �>��֡�O��ؑC~#y����:�7��Ɯ��x�˫�n�m��|b]l�j������0�p�u5f��$q�����c�?s5��aF���v��Q�ZEe�����qd�FM3�\�k�g��C�3

s7���8�y�0���N6���(|����y��\����߮�rR;����i���'0�P���k���;/0�n*�*�9�������Wf���X�\/N*�"3�Q`�n1ݽ��;{2��M�����u!5�w �������z��DKA2�￴�%�$.jf ��?TQ_Uh�>,;���a��8Lpx�_ӣp��]t��D����L�6�ߔ;,V�p[[|�;p3zx:���@:ciFf��2�A�V�i���{3�Dg��Bi�����Úx��]�Xo�?H���5h(c�d�A����RDTg���J��Ŵ�@�؁��ǰ�����˕��
M2V�|J���	�+��/,���*�N�%���fal��fv� Blg�UQDI�Ddh�Ν ��衽��iD�,@!ℊl��+1��c�j���k��꥽9s]CAy��&�ye��r�Xa��c���w��-��\����tR�n�.�F����[�j!y�=Y&�T�=v��|ZZm�z�[�� �!��^dŪK��sk�\�]�#m�Ƃ��O��3����WB6�/8�e"ft���b����s�h���1�R�<���W �h�Q�/~=܅q�s�oɜ����nڊ��9�k���c��Kv��m����n	$��xP��؛1�{W�][w5o�
���� L���"T�23b�w���٧��:pZB��K��XA�����rĖ�V��	�E%���lw{{ڽ ����^9�<A�����l��PX�=��LM,��6�X���Q�fh�G������#�����&�!t?���wu�� �6���~�C��7<�LA�m��:�5�逞�v53z`�ؽ"��=��{<G�p"��X��ę.�T��ml�[����t�|,�GM��=������0���l3��e��Kxӣk�RO�>/f�����Z޷!����T5�c� ��G���M���L�ԩ�H�q%$��2|+{��4�a�\S����	Tf���<�������~��ٖe
ד�6�^��Y���G�'
�� Go��r�0�}N)�LL=��n�S�f/V��F��SB�������Lx��~�h�uy��Cah_C�]Z�H�d�W9KhuϷЉO�D�\��0�k�jD{(]��6rif{/�Y�E����s���I�"������pg��P� �]��������V���O�	Z�%qUH����ĵa�t��H��?&����z��cg�r�������j��w5d����)���R��մ|�N>o�O*�d�f�0���ք�L��e�����#N��9e��zT���!8�8���˵����t���:ɶ�i5
+#�u�b	G3@G�>Og�V��u&�8�W�p$%Q�J�����e�& �0-�t�Ò���9��TgN���g�=��_:ʷ+��7O�󾦎{������&4�aV�m��<P<�'e��:.�Gw'5��D�P
6��l�^51����y�`$�kt�.QH!�-��_��6]O���"A�]g��KҜ];*�(dsT\�����9
72��`AÓ�R����p��\��B�蒳��7l�}�ąBh�U���-�~ؒ�Q�����&A��a���Re�����sJc�𞘒�'9�؆�p����ѕ�J�7��v
-,оH딏�J��݂�X�ݳ��uxTA�R��'��+<g�m��46���i)�x��y��g�:�P�\;����VR�m�����(����D{�j�N���	��¹|���F�l5�%��M��J!�)���مf��r�V���zQ���ܑU��	ZYk'�=*�ҫ9�(��08��d9��=�Ӛa�ҥf�Ik`]Q��S���"��G�=�ݲ^V�F1ft�y�<F����,e��Lo���ra\RN�8��ս��.Ύ�`'`�P�l\�(��(�]&�s��2��0��{��>�s�u��-��3���%?�����L���<���ë)Xx�G��K�� L�!��ӈ�C���*�Ůˍ(s��j:p�3'k��K}8q�����;�e2�	�L��x�.�����]QMj�-70�-]���o�T����m�n��d��
����4b��~�n¹.͘�0vή~�W="&|RЏ�(��O+2�M*ͮVjp*ld�qj�n =o�z�[�Ʒḅy�Q)��
���:8�@�l�X;U��aN`(�~W���'2-]�Ye���n�Y��#��;���M	��O�0���L��CX՞�Y�.o��P�a�uM�S^��3�Ԙ���+Ov͙���Q��Cw�NT�-z��Rh�8�8�b���3]go�E ��|���1�|��Z�����!�] ��)s�S�ʟ�_;5J�a���c�f�{{�+㼴�]�6�c�*���Fo�7Gő�#�����*�$������J��}��a�ڮS@�� ��_����?j�
�����(��+���8]g�o�Ʊ���Z�`�eN;C�uk8�7���G���\CDD�>�冀� ʻ��+�s�ei���۳�)��#��m������ �h9��W�_壞�YF�h �SC���W��8���[�ɩ��e�\�»ڛ��r���R��؝��$�(����&��U���- Ra�ȍs���ћ.��o�T]��t����/\��i?��A��Mο-?��n;����.Uȶr��jh+�s���X:p��W=�Rp�L�g���J���Y�e�1�ܹh;�8hi����q\?Z5�`Rwx��'�ws3=���|v`�К���n-�܃�)��|���un^�1��k�(|3�	���Ϝt��;{���^w���h�W5&�L�F�3�l5�kU�^��Hb�@ar?5n�뛚�����3�9 }7r�r�.�wt�%�GF8o���Mx�E�:ߌ��HRaI��R�C�Oy�x9� ����o	w�(6-����i���I�������eXK�6,8��%$�Kpw����N���Kp	�����ۻ�y����73��W��NwWu�-k��n��r=���W#�dXz,<>w��-+���-֚����а��8[��'v�����t�>�#0�}�� ���2m�����=�Au�'�g0ؒb�Q�cj�{k���kv����/�@�C9�geM�it?��+��6mA�>��G���R}�q֏_��������V>(���tśP+#�e��<xѽ��ePƶ���f�I�VK�c���9�!7��8��W�=P:�#�n����P&qߖu�\�����E��Á9+��wQ�q|xx�T~���hߑy���/7�'�@Q.���W�PAT�X��.r��)q'\Wp�B%r�����L�����]@E	�����h�w��m�|aP�gNM�1���sIx@@�uG��*otr r����B�l��A�$w�cژ��e�q#�&�����Gt8�s���I��j�J=������*#,������o;~p�m��yK�Eyԣ�6: @E�]5�J?:��r|�Eae���k��N�uҴU��� �?ƪz��"�n��u[��Sx2|�;A��i���DP��_Xh0Y%Ń��{1v��$�/t�$&����:�hX��;M��'���@�9 (�^Ñ'�a �jه��`2�"�_N�4>�)�%x�~I�e|�>>���C�SMJE�]2�Vc���a `��J�3��Y"f>`�lk�p�G-
ݻm�BX����I�D*�U��_/g���~(�ߵ:98$� ���g�Hg��d�h�F�L|���T:4��N���8~����ŧ���t��D=��@V�ը�ͅ�+�E��B?+U����K��*��؀�Ǜ+�5tI��eк�
|=�ÿ����:,��S�Z�D�m�Y�L���DX���:a˖�����Dn2a�C�L��!=y��(\�n�zR�\k�v��itG� E�� �	k�v6n�[v����Yq�l��1��zה���Y�#�F�}�2����˖YOq��&ג�;�����VtВ���:͊b1[�ʓC�=�����"�����/bү4h��[��j0��I���,�
$���lY{�AL�t��[PB9o7+G�a�mb1_��w���Y�F�5#��^AOW�C�R�i+���#T�sj����Qq"T�X�˞���P��3aꌺ�{����wI�`�4�'X:�`3�cqz��	��'O�
�n������Q�硭�c�/-�T��wbL�1���y[E	�K�v<�Lu����5iz�,)�Ŧ��O��� _ǯ��*v{��ȹy��
b�f��^K����>�W��C��k�"Ր�퐷YgE�4��{��A��L�ۄ�=4�ݫ�����Vr�k��`��gV���W���[��)���۱�HM�]J ��.�H�d$��6a���4��y��� y��}�I����˂hs6������ĥĄ�&	��̦�'G�v/7�Z���WfD��l{���>�}�}mҙߪ
E�`�w�� ��1�ߔ
���ʄc˓�/ 2�o�@������ˑl2yPFv�6��x��ɖ�A�hW��+�IUrԔ;_w�O��'�̀��lp�TU��6�ik8u��@���cy[l��9��#n0�M"�i�����~���7K��S�|秃N��{��:}Cg�Y^fz���DԦ�J��b[�2�KW�0���6�0�Sᣟ�-�M\�Zd�o��|�l����T�g��6�����.�N�o8^�.�{<ZyC��}�܊��5�~̘�2����Fx5vR��gR<uCmײ'sP=\��c7}���[CK���f���vI�c����W��-�� �!~����t�����G�R���a	(���=�]YT��[j	��\շnIw���ݺW�`�n�����ybU�(���h�HȪ�m&��<�ʹ�O��JϽ�_�~X���R�15�~�מ��=����c�O��D���FT�J�ex0QJ�`Ϫs��[�����{G�Y�eSX<{��u[1(q�1�t��z�d�|�ṳ���ږi;�Y��ב��߫���fý���2M�~j��܎OUyp�^IUW���D��g\��t���?��CDL���/�1[��K�ξ.�&:m��{BL~��7%��u�@X�nj����􍸛�*	fu�h0I�s�m�0�� tD��M�ۋi�G���];��Vz<�]O m[��Eհ���ۼ$�A?y�F�h����K�A~�!�)*'_�ҁ\��K�YPt]���71!,������4k��S��}�B�~t+U����˼il��C�j:_�ܠ���q�]G�U%�FVW�P�o�Q`��ـ�H�,B*xZfV���2S[]O�y<��2�x颟 �����~Z��Yw�p3��Z����ģ�+U�	̵�+�������vzj�ӥ�'����7�f�%b����-AV��t�2'�d�t�ɋF�:��YⲺQL�c0��:��uq$Z����˴��^L�K�
͠EU�m� ���Nӻ�:7�',�/�Z�ڴ9�g�9����c�K�-fh�Oǐ
�7��e����"��VL���C���(<y�sy;�be����-�09��K3K.�����l�F�d������"��U�j��m�V�][�^�����[��ݯ��6/�G��x�y	��Z5�T��B������@w���޸�V߹W���@7�%�k�8]�W�6h��Fi�^:WW�Թ�J"C ϙ�h�t��>XL�4Þ��6��ws�uw�n?п�?�q���iE_��$*�L<<�h�˲2�C�6x~�P7ف�.[�F�|-u=;;��-�+d�A�3B�2����^�V�j{�89k���Hv��:����of�[ߴb��/f$z�����,&�9�cġ	
]�5=��

¨/}�i�UƳ煭=pa�U��v��������,����?�wY{�t��h_|b��[�}־�$�PBUJ�F�������>���t�P��r:���}[~?��J�y�92�s���3���A�P!E�GX?g�|����DF��UG9̀��+�8BY4+����f������AW7l��Nv�J圫����p(�Ϥqy#�<�g\����]=Z��px�n?ߥ���5hI��lbWi��n� �̃6d���ބC�5P^���[��V����g#>	���z����d2ۮM�h�Z;@E@�__�lתҎ�G�&�@͎_�}��`V5����.�:D:fL�-=����;�����b�!$����?5IT���U'�=��oh/�5s��S��{���]�6�\��}��MGK�kX-r6D��/���3���B)^�Q3�|��/P(�i�xw����Q�E��1��y��ը%kgQ��[5ʙ�4�.K��_0�6�xP�'t���nG�R@����E��۞�W��.Ǻ~��P��E�2QkV��|�5_��r�"j	r>>�LY<�0�i���~EG�h��9I�oi^r�>�?�Ƚ���b
|j4�)�p����?�J����N�}rǁ+23R|�`��=
��q)������u��R���f/�ω�0��8P�S̎����܇���~=��<%ᨃ���w)M����ۘ\5�1��(s1E�����/��c,�|a���Zx��h�K�H/ s��[�V-���(J���7rH%b�c�}%�g�i����`��n'5}���H�ř3��@s̼�/F�wp#��h�Î����G�l	���&�Cj
_����/|��v��?|	�ì���?��g�H�,'��t��,�5�kŞ{�H��c���q]Ƴd�W}�x^q�B8��ᛉ�m5�Kf�X4��HZ�%�����m���[�R�8����z�R�z�)�R��v�(UP` T��.''���Rt�����]��,$��¢��������sJ��Bs`_^-/N�
��vȽk��K�"�u@�;w��b�ph�ۧ���Ok�>��3����V���QJ�ʮ\��9������D�'��YW����Z��X!��3�mS�����w3�4��N\���-�Mglm�ډ�8�{�L��'r�]3�}�$	���D�Eӝ����%���[ь�}������� ����e���@+ ��To������olȄ�a�d�/��%�bf+��z �͕�g���:��VA�X���cyYܻ�3����e������5~&�G�(T,�8|���ȅ�<�(���:���x4:q�J�g�+#���4��}�D¦�����:���B:��8]�oͥvt�Q�0��V������^qpF���N)�<dA��mioId�(?� �n�y��ː�u�\�>G�����ͣ�U�û�����_���ΛC�z�܄=��BNN�7��9���ež8ޞ������1.R���P���*&z��15�Ӎ\E�'�=zsPw��fB���Ug���P��b�xP����a��
�~��B,�n���M\�:�'�w����>�m���5��N  �Į��I�\�O�����a��Z������z�!Bl%��^h}xŔ��������(�W��ݢ�a;�T���I��u?��&���+M#�	ԩɹy�8���ݧ�Y�/�WT�۪�@��YF�S��T�߶���]Z�a�\�ܼ7��9��f�5$Į��� �/Do�5�{wc�_:�9�'J�i��vJ���)$���d�T����Ӆ�f+.�8&���]��>�u����TY�\�o�7Z�LImï����z&�pL�����Kk�t������{P]^%E�޿��m��f���w�o�[�Ѻ�:*�b�Y���"B"���0_�]47'܃Ѳ����r%��T��h#�vY�v�=�KE��'����@�.���L��o�� E�!����;������h���p�c�^����#ӯ�fg�f7g�A�xŌ�R�;�T�����7*�W�6��G�xo^6q�)-��{�@wۺ-4�*w����^�7�Ω�.k
��$�����>�(|�/���$�'&�m��â:�J5�#�� �_c�:Y#���:J"p���)�u�rZ�*n@�?����޼��h(+�}�F��EF��c���XihkX=��4t��?à5���4�nT!r Z=$rd��c�<�>		�o�����mO�#5:�{�|=��gJ2�.����%�o��o�����IsV=�B�~��<4�5��]f6���W���n��(���o�+`�Fs�@b��J���˂l�"����	o��]�G��k�[Oy���Ob!��f���4I��L���I4\�6-H���L�?�M�2� ��]5sk�p��f�ݦ�Gb��� �LX��ĭ*o����]���]YwS'_��M�c���޲�F
��k� pFK�r�/$Z�[�];Y�gV:Ou���@q1a hϵ&�ÍI*k�*)�0��YGO�Uj5����6+^�س������r�+�����b��O�|�{#��L3���bX,�'��3y��j+�oh%�3�?��0�� ύ�N(E�8��
5���wz4���,��,�����s�$q���=�3���=w�@0�Р�]����=��j��RLqjaO�s�x��t��=������٧�Ks����eO,19{�A����a"��#hх�s�>��������iyn�K��-�pN�]�T�RG���= \?��C�}���0͊�<T^�G��4U��t�{嫇��_�"���)*��񅙇V���"+��>ee�fy�&�Z,oYh���i!wN��F;3[�W�D7��ʹ�a�Є��`I��{��2�'��D�o��W��'WoA�̊�R7��C�/L��A(+��夆�/goZ����p�����K0��CXb�_+�g�-��,PH$Hr ��Y{�L!#�X�\���m���7��<R�l�Fn�F�T>/Z'�N�M� �b�KHHL&�#`\�����i�=�O����@�	{*�?�C��<���M}(ğw:T*?c�m�%���_���)R�g_���;0Ռ��4�T2���W�|G`�[[t���(@A��Λ�����s���@��a����l��N��a��8��8<Q��i��E|�,!=dԏ����xj�&u�2��A�	�����۫�yz,ߙ��p�8%46oD�r�RS$
�h�����F�"���ƾ5�{���z�����N{��M�*\��j����@�
UdK���hS(��?�������w���Cx/�現��)�������Ј�&*6JUr���8׮�/��):�Y�����W5W�|d���G9��G�-��q,��Ti��q�r�[��vJ������,�Hhx�<{l˘r7��6;Q؏2�FX�P��~���RseP�u������JAhp�q��_)�2Ę��$���FqtY������`2K��o��%����-�rv�7���Ί�ф�3턉���ᢠ̛�%hŤ
)�9�����I�0��!���ԃ);���㖤&2�5kv��w?�r�c�q�}!���6-Դ�؞�:[��>��N�GE���w>k�{Ey\+����'�-��`�X�1˵�`�p|rXQ�4bn��[q� ���O\�t��z_�T��F�=gu]�N2�D�܌����x.Cz��.@�R�v���8��w�J�ʋ�7iQ�~3��PN�8>>�"����YmԱ��:<<���U�n�1<ě���|A��$���*&���(v�<`��	;��=��E�۩�0�{����[��\^%�xC"8�+���~w�Ȣ��׊���f
��N� ���c�6�I�'�_�����SC
����Y�3�q�IӦ���i���>,�P1���+�1�4}���7��4NԸ�Łؗ�8CbE6U��(d0jcG�i`�թ�\��0��A�<M���0��;�]��1�W?�5:a�nx��\��+���qT؀@�(��tPj�dk�t���xF�ĵ�����.�^��煩�GE�;ez�о�}�u]Ӽ�����IR��ϑ����ײ�7�)ɣ�6]�^8Mj�+ɓ���J���,�#�:t�Ap;��vT{���~�ʢ�ݽ���z���_��~p;Q
��*�7�4d���'s`�-l��'<��*�������R�
��ح��;k�՝���\�F� �/S��m�ll �iD�M�h��B��!T��8��U��W�Jg�h:�u���t����,��@琣V1��j���׫w�Js�ph���>���f��{��o|���y~��&Y�F��lmkk�yϼ����d�x��)�������i�m�Tdld3�!醌%���t��g�;��B�H!�����,��7���)���]k�����B��Nh��Yϯ����|�`,�5���q�Ύ�u>�[=���o�Fw䢨��1�g�����E1�W�+n@�M���0�	��f<T�U��������N���^Z�3�
�?p���k{�=��UIv���3���b���|Y�^�q{�(cE�C�^ ���z���E		x�5�V(�^Q;�J��������x���������&�%��eb�|�_���/x����kԛl��W�l������1l�E"���rG8�d�w�~K�L���:��u�]6�%cҨ�A��}�Phf�-ZnCd�sx�O�U?Z��:��c}$r|ܿ�V_#��q9xCuR8E���"�7H�j���lE��S�퐩��騼� �%�]��!:�X���X�˔��І�����'>Eb�8|�Al'�Ā���ԑ�j�_�2)�S��^Q�f���>��v}�!	pF�paQr96��m���V�Rg��x�x:���b��;�_��7ԙ�\+��,)�+��~_�`۫�"���dWH�qPu�Ο�4��(3[��K5\�/gt�������̮j�wRM0H��nO9 Imt��[�Wԋ
SPZ�]�t�6��H�>�n�%_ ���������-w��/�~�1�>�YI���ǬTK���ʫߤsW�Lq�j�x�l>�@d6�C=�E�5�~�8�`,LO�G%h�}�g�(ˣ��Y����{�s�p	�����l��}�a��B}��샥�9�-����_���4�L�?(����	\4�P�f��/��e�V�O���f�Es��-;���d5�@���tPmk��~�˵�:�c�6&�q����o�E{m�Z�=q3��0�`�rL�]A�^_����#�0Xo�D�fj@C�Zl'�H�^�
��u� l�e��S�h�[>cӴ�Ԉ�b�B���@�bCx���z�0��\�mmMf!��<	#�?�a�D���P���)��R-ri?���3����
�H�~�B{����H86��{C�D zڴ�fu������-��5�	�_�a�+����c��t�9�h"uzvk��	܊pn��V3N�j��9�2A����j�E����	�WY��SqP�����A\�����^���N
GI,^�'|�tOpokx[՝�[���ٰ�#�.`&���q��J�,�(�,r��+��<��Q�A���ݑ\tS�Q�^r���B���z���M�U����
���`��Q��1�i�o�ZY�AQ��賰�亇UQ�[���1l���F�r�Dpz���އϯ��D�gl9�a�b��o�M�Nm.�{:�8P�ۋ��%��w�hmn�)*I�œ�⮆��5��n(�Ј �L�u<�����:C^3U��]�$�=8�7�����ߢ����ΧP=�8��wo�N��a�?k�hs�z�u��@W���^�r[|��HLpJ�yr����s�5N{�3N����n$Q�_Ą8PCɡ {�n��a��҆p��B�I(�%���PP�܄��Á�����q�L�3,��$���8�5���!��v�bѫ�R��%c�.�;_��/�;3�҉�iU�t?���:;DyJ7�ƌ?��t/�eP�*��6��������6*e'�e��G�>~���DP}B���E��y��vE���"�O� ���Yw?�����"�i�Hz�1 c^�<i�ߩ��8qp��U/7o9T��H��A7(�o&>u�R�>H���kf�TC<,�	{�]����=+!��,?">�m�`'�T�j��w���e|]����0_�������'�,y9O6�ƌ����˧/2g�5"��oߓ�~c���rQ����/���=
]3^ҁ�`����?�II�0.�VzLw\Fl�'!)N2x�o��)y����+<8Z�퓘�T�۰��m�X�J=~Vpq��W�������,�s���;�٣ߤQ1��E�C��Ҙ髉��Ѯ�m�"F|+��B7�,�tq��;^?�O��{�~�� 1@�ai�(���"��s�^�qŪ2� e���mS�,�'�g�T�������Ng���� ���cԖ`�ۑ ;��Y��u{�[š���9�SA��#���;�[r>w!�p+
� �{��x��-騴����-�~'+EW���|��_�}:N쩁n��M3���W��9��]0c��;�������-"���&f�f�`�8O,����P�O��	2��B&eg������c^$�$L��?�n7��P9�v�Ѽ�$^ ���B��T+�@j�����Z����C<����O�(��^@���>5�a�~�Vd��6P8_�CR�q���4~۴%,9�ء�*hkF��NqHٞcT\{j����<mX��?"9߾EɚΡW�VU�s����9ڄ��k�v��T��T�9{���	.h���}^�k�wv�m�Y�g�r����bNZ�<�0�bl�(�;;{�s�	1���f�E�C�]�:#��PHv*�~�=0����j)�+J+�P�U^��@ğ���Je�߻�͟�"��c�H�H��1}��y=8muI�r�����Sj�K[�1�N�ٴHR�E�-�t7ݳˬg锑I�G@��$= ��o�qsV��g�������&�؟���}�v[�%�*P�'�myO&wX��}�uH�F���X����w�Ӝb �tB��J��5:�]�J뼰��hH4�$��퇰�Z4�~K-_��N��������O�{��PIk����"��ʧ�]���dH����_����[~p<��ϳA���i���v��Ѿd�9�-�y��L^��z��q��d��A����6����he2֞~�����$��J�����Zb���!oЈ���f:��9�`x����H)�-�A�hF~?��m���2zt�'��4����N�M�p���|..i����f[e�@Ց�Զ`���7����(�)��J'�]z>��L�'��M9t�C��9:N��a�����;��\��zH:��%m�h�r�n=�Ϧ�>"�L���LΫ���;�pߴ>+n��L,T�4n��H"��aA�L9S-\C�����*�vp����/^�
�ˉD#����AizA�
���B�C��F���4�%��H��������M_x�}d0V�NG}KK{�a�|�0�O:sdHB"z�0�]4���;������EF�ґo!�%Q2��2��7�q�ժ��"���Pl��C��
��B���-`�aW{�\i�bg�q��s��kG�^�$܀mY�.`�Wn0��P��n�~�:��w���i�!��;�PO�����5`WK
c2����馩�ܢ�P7 �a����םL8�9�>�g=��w���?v�L����=������^|s]#8��m)*?�kk��n�]�,�� �9*���7<�UǍ�Qg��aŽ��o:=�RƦe �t�\ɲ�Ʉ��7-w#\�|#M\�[ ��g��c��|	����b�# ��~}�9���<��J���k �/�z{yX�h��
�2B�p�`��?��y��0�&iz� �8�c��4�(sVH��4Vpެ
�X�x�6`����,��+��������}�z�� � ��uF���� a�G���!�.�h��x��oz݁k5����5j�Т��ھ���&R�>>������Z1T���D>Q�,���b²V���^�������ɵ���p�Y���<
��˜J��&L���G�E���MqG~ge���C9�oZ�F8�V��3��#K�g��������#S��v.y{�/y�5���	��<Ll˦`5oi��c�����bf����\,�/㏵"�2���{�����iZ�:�X'�p��nd��@ҕ�J�m���u����[d0rث�EÝ��"����j��h�΄�������I���@��:w��$�T�0l	q���OV$�SW�_���T_�(��|\�'��H�������{3�v�c%y�x�SN̥�����y�oe����ʩ�;<W@�(
�l�Zkб{ǜWev�4����Ԣ[���������IR"�>���P|���J�Lv�{����%�K��������۸�<y��+���P�B�ud�}��μ"x�5}�ѠT��T��&{�W->���UK��(,X�h���kI'�d�!��1�8<-h+�J��jU	��zY֛.=�+0����@�Bx})>[�ͣ��Jo�����B�zߐM�3�D���сfa���]
+��<��SkQ����:��U��>�6�l��-�\8���~e�i;��#�<F����.o6R��>b*��"b���Z&�vCh�qD��H��d�R_�3G?��_fLW�u�#1�yx_0b�Z!/������o������9@C�,CAJ��`��$�5��e�R�=�7����gM��E���s�|]�;4�t��t����Q!���u6{!%�/���ܹ,����{,�ע�/=�JQ\�B����C�Ih?���$Z���=�QoR��d� A54=��]K���ZE&T�� ð7��5���e��Ɔ_�Q� x�^fC�B*醶:�a; E�ͮ��*�2���lgJ@�]�~�G�>�����e����TPi��V�9L3�&s?	-�ś�� e����qR��\��m��W,�a�X� ֪9����Pӧh��Aw"1-�1K.|�u�8�>��V�H%��,��kbe\��
~fў�	���O�;���I:$T]�[��<���uq��;�"��R���K��%���Z��`�:�b'fR���)a�]�4���A�D9w=K26�R�{y؋�MC�?�M�ᕿ�����}���y�>��h:a��_����t�ބ��[�u:�Zy�'�#\l��Їy�����Z���hG3t{�O;�Q��t)���4C)�S�����������d���)��J��|�[��@�|�5_�i���<��q�Ky,�؄Hou�fP}G�2��Փ��s=�lCz�ߟZ�k����2w>'m1T�cۉs�s�Ň2�Ǫr�V�K�*���1s���-\��y�<~z�g�a���U�;��������4��a������ic�ܮ>�P͝le�%v�{���>�P���6�r�hD��{q��n�U~���	@�:P�|�3P4����]���3MY���<���|]��cI�����0ts���58 p�g<AJ�"P�?OzKf�fKRf��;~:\���e{�9�_M�ϟev\r�ݏ�Q��Z[���uĝ��g;+輻���H>��{\�2��	]�w�|F��Q�ŵ{����7� ���f�pЬ_��֧O�Y'9m7�]��m���f���r��`���in�ϳ�Jb~s ��V�
NI ���+�4t��]�>��v��$��p�{>��|p���{;9�h�\� m�;�;�ha�w/��c�6t������E�z2��hɯ�Gx9��=\� � ��V�NnQXmj�ɖ�[�
��c����
�����oU:���_��ڮr9��� �E����B���U��)8�t��0��k�""I	W˧4�<�Y�/m��O8,�|-pLJЍ`�7�X�q���N?/{gQ�����,�C��4P [%@l���	�9cu�;_��%!iސI4�ǀM��Aޡ�g��c1��O3%��$�S�8"���c�����i�\'��{e1E�+j ee���?�Q�]�k��s&窈3����6^�L�ǧr��Б2A\�S�6���k�Ŀq��RG:&~�L���S!�ѩ��͝H�L��_�
@C��8&���Z;8��,�8ӏ�D*Ĉ:d�-y}�i�;	p�Y����i�9qLS�~N�L/�=��1���PBMW�sv����F�l�F�j��ʤ���2=�Ѻ���ޮa�M�o(N2$e{�e3�%���
��#�{7�4-�}��["�Ug�\�g�W������(j�Y|w�}q��'*� ����:{�G��$�MFw:Y	&��%������2#������S�5��9~	P�% <��a��H$ʸf(��W��E�p\-���R��Y��`�e��G^�Z�N����YqQ�w�h�/  w�u��8�>��z���݉�T�����;�ڟG�޿�a��g�-P�������M��o>B0�wգ�W��~,��}N{�&i(�Vp�� ho׾fN�T7Z�0�O2]Єu�ٻ/�U72Qh���Jq5�؅��;Jl�(�����e�� S�B�������+>��X��֟'Q��H�H�t�O�O%���!�@�� |_4���L�Ƭ�\%�Ň����`�x]H�RY��(�fo'Q��W9N˩��E���F ��� �|Zr{�ܰ��VG���Ɛv�\!�6S�k�Ѕ���	Vw�ӑ��J��Gћ�L�j:^%d�B�jh8���G��r���a�՜��Tc[
]��\A��+��\�m=e$�SWtM�Ƣӵp�{�\��d�|�,�l�1я�cQ7���hd*��}\("�\[���0&���>����b���n8$��h�}�R���%"����GI�9'�p�wb��t+�w����]���IVO���TLo��eRz�2%�om`Ŀ*3���L��,��+�h8=
�VZ���o�`��|�-R�+�/���� ���s��N~�x�8]�w=�d_V��V�B��/����c6�Ys��v����0����
�`��
r�m:|�M_�[�-�X���T���+���I���\�ί?���V^�i+jэ8����u:0�Auc��1�ty�X �p ���U�jz8�x�b�Pu9�жu���Ԕ���єi�;[y9�,R(ƴ���P_�v|%0l�C6Ou��ih/' �͜7-�B�C��}Jo�����$��(��(Թ������x[`%�q��a4����y$2�I4�(�͚�]L~T�	���+u~����_i�N��X���.8�t8Nv�rӮ����V����D��%�G談�B��/i-�Q�m��n�N1�G����^5P3� ��3��`���z��g��!�$nE��k@�h��?�:\E����Ԫ��ǉ+f[��[��3Yl��m��M���/�낳����*�4B�LuJZ�qm�`Qo�t
Z�*I�z�l�C�S��{��C7�Cqx��t�a�&* ��>���v��	�csc!ć���s���D�������<�r�W�Y��,\ơ6տ��@In�?Ԅx>7v�B�U�~�{	������*T��S�~7���i��4�"�:K��}��N��|]x��+2�D���B�u�n9�[��󓖬���3���Ӛ+���V��a��x���6(�9IT��
��0�x5�P=�r�
��yb\�ҞK���as�t8��+���i%�?�:���R`8iѶ��'p	��B��;��
u���d��+f�!��u��Ҷ�NX@��3��5_�ް��R���li�/�M�@�����2*
N#ۢ���-	���'|e�ҷ#���[�K�m�^Ü��"��F�Ճ�]���uؕM
�����Fd�E�u���}�3�����>���`;BҜS��V]�}Ft�:���zd��	;�2�X����`����;�O��_����(�*&�b��e���`04�z�kƹ���{dnXz9ag��Z���	����h��k^�� ���]x�Ľon�E3K�ל���6��f�?���J %9�PH2C�<���y�G����\���k�t�芨��D�E%����^�2�#�8�I)�4�p7n�'V���7��B~�2�#���D��S��t~m��l5:�;�7k��L�4��k���wp����?�_��>��)qQɺ�;��+�b��&i�R��e.f;�%o��(I>|��Hks^��Lj�!H��0G���T��7��>k��dD$�ܚ���/�a�'?-uQ��V�q7�]tn�t\�hO����`\y4� �Ԕ� ��(���-�Z/�79�b��Fή*�\¯���=Z�����y�ѥ�"�5�T���d��Y	���g3�M8����-�n=�Q;w]�����f��7S�N��v�yi�����m��5hk�
����2Pu�,h��@V�qk����;$�5E�l�쫿 b�[ƾ�LG&P�~�2�C�Чs��C�:|�x�a���{�^����};(�� ��Xe��Q\a���H}=�f6<����&��]�(�&��T�n�J���撆R�W,�R˾m� �m�f���8\H�lP<&�J���^�E�hf)�>jt7*�a:�ԭ��w�_�_\��G�n�%�>y�.�*�=2��2
ڵ���v�'�[EK��i"��c�V�4�^�v�����߮$���y�"�U�9ĉ>!�����tVq�}c��0
��m�A���v���BU@>��<�5Q�N�ya����w�]P["g��c�ͯ�q�b��D�y�jSk����;�+����ߺ��QutCo9*yH_�U��UMn����mn��J��"��/H���S���Eo�l���0jh�9
>�gb��)��Y��|̄ku�pe��/:a��<F�
��g�~Ӟ�$@�(aX]���,{�_0B�������>N���$tR���҂��5[��i��C8\	��<�^�r�s�a�r?|�^��f����nⵐ�M� ���M�F'T�&�d�A+{2
^ן�t�<��S�u��>2s�2��+�\�������l;�w(��$_����}} =XR^�7nk�A��7��ᝃu�m+���LL��Fg�K��B�&zk\�+����|���Ptx�*ԛ��e��Vo��m�8�Z܁�f.�:�朴�?@)�*,_�9b�������\1w�cW1l���`t����fn�=�Q	��Z�c��7��ʫ^O��^�9���I
6Cn���-x��C��(��W�\D#?ꂤO�v}���'�ݜ���!yj�x�&�G��Z��&����黊����]���L>�gܨ1�2�
v#oj�!O�V�U��q�sh"���/(\�7�ڭ'E#b�HI�"�ŕ�T�F�s�x6�Y%������%n�┹p�K�'f���}��@
s������O�+����+��6
�屉Q�Ŏo���a�0�|�\e��6V����ף�����M��ڦf��}N��5.@��;��#3���&Gk���K}Ul7�����t'u)�P�4�M�g�B�W�VA�o.S�%`K��{��.6���a\0|ƾ�n˵!�]L+[��fpǣ@(�j�m��::9�Ԯb�V��}xUx�.�A. N�����u�E��9���UZ�{�6v��:!r�R���{��C��U��J�b��<'��Aiz��[�(�}�Y-VC��N�?����;�J���Ĳ?BFq� ���u�B���i��/~��d^��&`�Y�Z[�K��^ ��Q�v�q��T'[S+�Oo�(wÖɓٷ<Ŋi�e�ͩ��)N� ��"��'ۛ�Q;y���kW��b�-�Ŀ�pp��ާ�G��¥S������v){���eT`�5� � �% ��� ��w��[����Bpwi��h�����~�ٙ��6��z��[ϭ*���g�	C���:	?QV/�Q,In�.��ϵ�.�����͵ͼ�p%^�L��A�p�S�PŘB���焽�E�o��W���p�8G���Z�eRx-�J�UC���}�
l��3k���d�����M�:����)
�?�Ұ&C}�WKR����~۹��r�0n�W� �\؂��nzG�cx�aid&C%�'v[�2�\ei�$2�0�A]��;E�[���!b^��n^�0��aP����Gކ�h/�����6a���(�E*�K�Fl�b=N�z�y���&I��W���v����G/C�H���&�8҂dd�� jk�h��hJ��;�E�4��w�Q���I"G��Ƞ��û�6��z	� �:2�C�� ���k�E��A���lݾ�/�|���nK�Q(�:��%�ټB�,&���L�J8��>�?� *RPpXJ<��sG~4��:�Yb��ᙧ����.�*뎎M��$�<,���|8�u(�>s��`?��<d���r�&Rm<��W%�?�>*��}b)�G4�S��\e6��g�{�O���-+]咤�.����������c�Y�=�����S̯���,Lw�8f�T~J9T�{��׊L�s��ë�_(��zE�1�iD�1����T֐��\3i�%��o�CIA�G�E]no�����h����:��� 2���[w?�����5������]1wha|2�'v����r��k��q6�/w�{R��a�f-C4��'��$a(V��-�1�ܹl��E>�AN*������.Q�f��U�U����	%9��2�AG�7�11Q�s��W�˚.O�f���>	o�� �y�~��A}���7E�Vy2mŵB���Z��ۢ�58�1	3`+��Y�����𴩓*s�[���y��2�lRB<��ʅ�B7����iuϫ�������OG͵b�|�T(8R�_cz]�=�2�8�K�g �Qӊ��0�4��k�<6$���`!n�U�$H��{���{�b��3��b��Q��T"���%�B��j$�� �Nj�F��C4�� 4��A�.�f˛n���d�|{G*��sO�A�-Έ��Y�)rx�k��P��>L|�+P.~�!�>�*u�*Z�������.?r�[(q����.�H�k�	3c��`R�ۜĶ�7���מC:�ޑ�B	ܶs�א�R�u�!5	v�(�O(q�%1ypې
(����Dv P�L�qJ���=�hq�y�5c%;�V���I��W�B��&Ƥ��q�c^5�`��n"vZ=d�~�Rf���ߘr܅�k��%_a�+7�����$.����c�ȩx��|�Ρ�g��u�Kn�-駔)���QK+�s��yñy,��Q��G�K;��qO��v|R8r�	>Q^���V9CxZ$6�K7�!���/�����Q��	��Q��z��X;'c���OG��h������kY���!C�u���e���~"�x/��^C�Q!~��1�A�#fK�D0���+�k�*.��jT�rpT��4�BS��v��%�m�J��3�f���KT,�)���j	�q=�1��6�=rLjD�P:18�!ysdKפ"��R�*�fjT�TG��*��2[x�ʞSv5��yߛ��,IU�~"9��,B@���d� Ŭ!�k����k|�2��x��,��wХ�O{�3��G) �^�`k���\��`ȿB�:�6�)s��� 4)� %[�·��d\���j猃�q�J�>MEƲ2�ɫ��'"��f
K�o����J���u�0��N�.�x�Z�o�rm��M.�Pu-���L���������v]2¡ޚ��o /o7(5�6D2�px�#ױX�e�M����`m��~wp>D�O3�� Ш�ZӔ�p�S2���m�qJ�ڕ���5��5��_���f��ґI^�%�N7ۓ{�ߐT��!S <m�N�[!I��\��q�R���2a����@n��i���B�s�B�|3斔�o|K��`=˅%��>�>��U�6��ߟ�H�l�h�V�n|�F�X�:�v�<j��aj�
�Ʊ@iv��i['�ޮ�13E������,t�]��JG��N�f��)Ĭ�i����>�ʟ7���:N������:"'�s��R�����J0%��%w���S��"�����B�8)���Fq`���K�-?�ܫ�{Ӿ���D�	�\>EK���@&L۝�\-�y�I�}��m5�<q:�F,.�/�W�Yh�Qަ�����ǀR[�^g�x
��"�v�k��d�?�~aR��&�����c۸X�i�@���2!��k�C9-g�F`������]�ĺ�S�?m��U�9�k�I����P�	�o�MjNU��>�$�v�l���ߖ�/4Aϯ䩲z������,�֖�(���P��d�%�Xg��/&���H��UlP�[:�Y!�
����?���~E��fl�78��cΔjҏ�H� �h���QL�.TF��a]� ��w?M�J�*�>h����<�ߋ����I-z�I�'� ^d+�z��]�1�
^X�h�+Ť�������!�� �	�8g��K����Z9���fm��F���(
ޣ.�^����k��7��O*T�C�"�-;�W���@�E1����ƺ��c ���۠���q�MF�S�>���C5�m���F;������M�!�˵�����s`��/0�v�]�z�D���0m���L���*|CW�k��Q�b�8�x|�r~y�[���zht�vˀs�ީѬ���x�����%$��_�p���T)!D:F飞
�(�!�b`�$<v�?�i��{��x�(�\`?zÚ:1��}�X�{�}���!
�( +:�,�{答5��0��f���w������
�BC�	,�s��𩪷T4��S�;��"� � �"3Ϥ&��&JU�+T��HV[��9z�^��^�On�q���V��;���
��MF�0��`�R�z�(�?����E|B4��n���u�kv��I ��R�ǒ�ʞ������t�.��|�X�r���`�<��7'��u�o��/^�P�	��H�燝v=�/ͨ�7���@��ܦ��� i#.����(B�J���m+����N�B͎��(�b�1tW���1<��Z�0��Ow���:f^#��,+V���L�P�7�-�7�M��w�Ü����c��Bu}��.'uU�߷�����GW�����V�E�
1I�5��d�tAFe3��aYIY��*_��a��2�I����5�Yn
�V"'<L:��f<�*�f}<�8��)�KvXI�E���\#8�c���zg;T(D,�s�Ϯ�8g%n(r�0&�z��W���fd��B�I��S� ��-��KL.�W7 +T�R�q(N+Q��ˣp�<�]��J�ɼ�£�͊{���R�ψ��O��8��yk:�hc:_�X�1^'8��h�%T�`y�y�h(�ң��B���\O�}_𒬪�/)�爇���P߮yW���/��ss|�?�;�C�,]���ӧ��.+Q֓����xĬvO�É
�U��_I����j���e�mt�;e�7 ����QY�����U��������U����r�D=�����l�s.s��Sϣg��FE�/6&��IW����͑w�J�+H�m�V��)R�"v�u���.����U���oxd������y���ne�:\�:�5%KՏP䷸�D��B�wP4�)[O���r�W�:´ā�e�^�|�o�h�-c��D����/L�G���b���3�ޙ�V�4�9��_Two9c`��t3�_�4�uR�Mm�{�1uZܢ���n~����'t��z�2g�|T��d��:	"M)���km�����ch�֮�#��|���(��b���ʘ��r�XSI}�z��}�R�k5Vl��^x5�I|ܺ�pY�>�*�ެ'���h�2]H(��#���m�#�>���.�<���7�]}lxb�+s_x��́��
O���9k�D~����-��F�
�����ڣ��V��$�F��F����v���C#p������L�M5MwM�;)�F��-Nl#�<�Iǉ(l�k��u�_�0߼D죊8����VO�j/�Dhsk��J�S�R�g����K*�&�A�؛7�F��n��Z�+�6j�?�O���l|�!�-�[�H��6�NmR��\n�R�'|]o�UVB��6&�0=((Ĝ4�(��4�c�>ky�-����ꉽ�Q:�z�_�ݼo�y[??1���ima�f����'��z��RD���+�F��W��p3_V�H��_�8��f��wj"���<[�]�V�p���/���y9ρ�=���aC�F��<�s�Z���������7>�#K0b�T��t��`�,��l��{���W���f��"b_��F���W� �8Y�$5����.Qǘ�-�4�D���Yuܾf��D.�d�:۳��8]��z��k;�z�JR����y��HTH���kT��譁��	�<i�e8�o�&Ϲ�¬��Pg�?�O���1�>p�}���+�|�����hy#���ǭ�~prt��)�j��2�B�Gz�pM8��s� V.�El#9He�(��嬳��&�ó!��&Tz'S�"�[�-3��6qh[ZL�V��NN�_���89]���1������ȝhv~zzw�
�2E�:�Vt9��Ӛo���Wp�X�+V׼��L�v%Ҍ���c^T������V�=��U�ˤ�`�ޱT&R��_��}{�P�+c�r��*W7+�(�08��q��wxS6E-����Ĵ�8z���]zB��X�qJ�aL�d�A���	I����B>��j �����}���Uvi����St�����Z$G(B�i3�J����;�:���:�����Py�0��U���hg��5#���ӓ�(f"/��L����ftO����WoS�4�������*��-�(�έ笞����J�h�,�"Xg�7>Ӽb�]%pUu��Yt&b�쁆�u���:_��*F���Gy-���&VK �c�uA������Љ�AA�����?��'E�
���쀫��:Zԩ����b�ߚ,�ĳ(��oe>n<��yؔ>�}���RKh��%�/��m2��m>�G1�^@�
Q��>8���ļm�x*i@�"5aJ_���t�[���E�w���P�Tfr*�?������J��z�!��1"����qqyP|��D��cmZ�D�K<��wUy��"�`
� �=�r��B�P��Ԥl0f���*��2u����X�wX��}>h�U\&�1rݬ���G5w�~A����G�����>���N�҅���*l%Ł.�N�j�lE��:�
�|�պ����ٴ�����1_ac&�v���[;_�H�V�m��� 뼒A^U���pflf���Dv�h��:��o0�����xQt�h{��2�#�~��S��9c�?�-[n�X���b��\�EiW�`��1� ֢b}��l�s�&����G1�!����o����������Ɩ�6g�*�A�����v�����6��,�����o�}�]T��P48��u[$�%�>G>j��
�gD�$@�����s��o�(�P��em�J�Xo|5Rǣ9�_bG�c���3.2ϯ?�X�?�G�oȜ؞�{t�&7��l��\c����%M	�J{.R�[5��r������M�S�����mF��ͩ�x���q�v=����Z�kƮ�
7�u�*�����kg}o�ְ���!r��pPё��Z3��t������D����fMG*��ڞR)<��<�ۄ�勰ᝁ/`�T.Ұ)�[#&̠�V��C����h�l%�I��%�>#�/r�tj��NS�J�/�N�2W>u:ݽ!	u������cmj2�q�_���HvL쭈��ȯ��1����z+k���
:c�	pQ�8���C�X���c�����bBl^3��.`���,��>!f$��E�r"�ESFqQ8/A��9沜�M�)�FP�g~'%g����p��s��R	h<B���i�?=]�)�L�#��I�z4pvn�z��YX�� ��x���?I�\׵���.��6n� �
f�I��t��U��y�[F�k>��=�}~K��dxe��8���ם��_��7�n������8P���"K/4OTJ�11�������/�F��2M=,cj>$}��IY���s�sVW�I��V���QQ1 �q�!�/��ʔ?ښ0�~��m\m�r�t]�X	��j�i��y���S��k�4�p^��)��Yz�1z��iXF�Qo�c�������o��_�ot�۟:8���+c`XM�����/��Fl-��ak����o[�#���9�ߟ|��TC&����6�Lų����/ÀM}�ȑc����S��	\G\��-�M�I'*�==���'��
9����5������1�QOxN������/TF�̾�����̆�)�S�d��+Pb�����4���}�Mx�*���n�V�25"xH� ��m�y��WZ�By�h�	�G�l��w��Px�։�����s܉���
.?	�3�Q�J��Ʒ��J� H����=�2Q�����E�����җz��`޴Y�VG����Cө	y���Si�@��K�Ts0�Ķˤ�u���@�	Oj������7���8/2k7p��R.L��a3`H���F����6Q�I��:w��>�� ��$~�)��e(8#�8�7�/��������5L�O�5�0��ޜN�#s����S�놢8����?�'2�v�k�.YF��%��6M�h��2Wk=d��+��za���X<K$�\�+j>sv�����W����S���۩�b)������4���mk5��困�&=��
�y_��7\%�N���Ǳ|�X�
�k�
�T�r��#6W7S{��XP�"��<����ղ��}���Zr(7�K�>`:i�:�2�5�Ps�h�,��F�G�9`CO^�b\�3d���}���jt+j]�l�;�|�՞3m���+����:��	bLH� �g���sS�(�)W�.2x ���g��Oz0F����=��J�||��ч�a�q�=×�?��U��s�U���c'AP�.���4��Q�a�H�U59g9����\9���O�>�������mqGTG?~,�7���l���_�>�r���M.�ծ����?T���}�V2���X��v���K�M����TY6�7/��LJ���E�5��H<�\�D���E�7?k�"2�dDpG�^�2�t�+��\�m�aݺ�kgI�\z�����>خ2����և1��]:T���p]��_�rI�F��=5�Mőf+e=���\��C�e��&��ݭ4ٯ�Қ�߿���;����rU>93�[����V,����wJ苄q�o.�.6b�8�k�Z.Ё	���'r��8E��Z���e�V[W[��RD[�GG$��''��u3��=X�j�`���83����#���~��*�U�ԭ�� ܲ�����	��{��OB箣�3�kh�e�f��� �Y���������Yb+����n�N��Fݱz�A���@4��t�����r��z����g`phQ��L�#��+Ἔe*��3���^!�Z�W~���%x�4r�h�
f�F;�slQ�@�%�_D:r�m%֍�.��?�O:����۵3>�B)�5�O�ZAX�s=�����'\�"�K�pZ�ڟ =,Ui}��Ӵ����~�]��p݀���x[����f%I�x<�R�~
�t/�h\���i�8�d�s�K�����u`L�0� B�7i� _�D�u�C��J�o�� n�K��ޗN$m;��D���fZVh6�hrV�i����4DS�\�&���ʂ2W�GjBCB2ت�H^"�7�9a����2fr����������DAz��UI�|x�1�e��p>[�nܗw�~��
�����ΥϛO�]�V'䒽sRF�}�Ҵ�+KV�V����͆K):����/�O��W����ޝ�=S�Xc�K�s�u��-��s>�[�G�C������/����V�j�n(�}��kK&���LL�o#Ԅ�>��P�:ll�RKR>94�d�֌��'L�N�f�ƺ����TRQtK�l~�⪽7�l'�׊y��NDm4���h�t��&%�1LZ�SҾ���m2Gy���3(Vn)�5O�������3�I��q�����b����Ij���D�~�j�g'��4������� �T�rN��=" NJ�ing3��²�:@�]S��:/0(к�Y��z�aFk
̆�� ���i���}��hZ���`�����=׆���(���"�j��Q0��7o\���16!��������Y`�����Ko��r��j!̥s�����M��8�`��7�u�@�p���T�CWq�}'�`���^�L7

�[؄���<��ԎT�P&n��i��=j�|�M�����*�R�yT��k����cU���0%b��R�s��I�rK��������(+��⽯N�K�^��7�G��sAB���Ӕ(��Ae����8#H�������� e[!��Cm<�Ӯ��s�����'���3�<�8�i�Yʅ�?������o`�z�д��JOi��|�V�Uq|qI�VqS)/��mӓ���g�Wa�Ln Q���Hᩛ�~W������ �����/�-��a�~���yv����p�e���uB�p��]"]��>�B<���]���ݐ;)��ش]i�%ߩ�����2!U�&��ku�&m�.q��a7s��9h M���3�m3��k�a�?��b�>�ŋG
p*Q�v5�v��fM�@�şܓpX�\���<�A�&h^3��81�|Py� E�zhS�˻<���&!t��E�h	�U����P�=��	v/�c�{�1,���O���Q�����&��{�v��:P���>����&��ѓ�s�$/ў�P�K��J,.���ui��s]76Z�@īH4�xո�Ԣ�	qx@	
	1�/�j�`��� � P������~�mH%Mm�\?�1T�!����^��W3��^���""�{e��1���͵s~cs�_mw��,z����H��矒�^+�C�r
5�������6)A�g�!XJ݈/���Q~�~�S�@�y�]3W�d�*�����P;B�c��}�l�]���;�(��\��l���i0U)E	��f����7��Y���V[�Wk���JF��we�7�������zU�zC.�`����P<r=��M�<�r�f�{68)[�/����>���~�}ڹ:-��Yb`���3�ު)+Qf��$ч�q�iU7+�b��'���G>K�)R6����א�}+�y'���V{%)��	ŋ���Dd#9���x�?�]���t������4�}�?�:=��[w�s޼�U�.�k�|�"��8y����"km�l�7U�դ.I.i�yj��l�fj_�7�+��|���9���<��.�oBg���Փr�{&��$���ր�����h�H
2����>Kv3���Z�i�Wς�4�&^&��"�E��\i*��04ĝ����Sd�C�d0�]︧<
w���4�����u��g~���:��n *<��)s^��
,sP�tS��2�ǻ�Q�V|�=*�5�8���x��c�L�l�ٓ0Q�թlj��W�޶|��Ϧ�[�-���4�5;A*b��x;"o����)=��5?�����*�~\��Z�߀�;��w=1=|w��76 ;�`D�<
��v�F�g=�%Wo2!�}�N��RF��JwZ�9~� M�)z��7jo�X��k�}°�l]WPy�d�e#`Z��JF�0ۤ�{����jg8��Uń!0���f��?�hɲLS�p�lu���k|=�9tL����ڻ}m�=��>W�7���3a���ҵA`�CQ�il*OS��Y�D>�]ɞ�|�0�����Q<oބb�q���PQP~7X-���ܰw���iT�/�e�D=N�%�~Hc��(.^D�a�,ޫY)*�*��m�N�b�^����C�8��[?Q��-%CusUK-��}��mi���rs\k9G�"���9KHo�b�~ܰ`��'��q���F(���rC����}���Y['��mNH����/{�ޯ���S�-9/]G]K��2t�W�iw����9J�ŵ�ǆ���I����a�h>4�݂w%�h�{0��d/��r5���Hv� �3�1�!� �/�wM��
��<���iP��ǝ��n�������X�^�:Mك���c,�~��ථ���f��U1�2Nx�,�zU��,8������j��`50\������\}����<�ȁZw'��.�^{GOvM��3�E?�W�;�+\�uҧ�̲�[�&�rZ|��Nc���u�4e�j7�,O6�Q�~䤜��yu���y��<+W��Z�2��E���uY���D3�61��]b�>�K��;\V�����Q�{RP�B-�S1�!&�������9s�w���[K������}���s�U�q�Ps�R�L�5ok�m�ti���k����q)�h>�w�n:~;}�� �����I�~����5++��)NN�������m!��O.v��˼T�'���J��-�7�&��(?���J�eQу�~�j���ڛ��ƫs�� �Z�H�;.�I#�)��q�h+P�GEC�C���9�'����^c�u�Z���Mb%	�]���(}hbz���)��6�h�׵t��[<XB��MB�X 9l*;�Yҗ�g��t+��k"��Ч�����#H,п���3��T�Rm����L�e
�@�i�'|���K��������U?�F��͞~W[�X��Z�>��O%"��k "�6)�˙.y��}c^+�S,ɒ1�@̮��L��(�:��[�>ܵ�'�Z��U�ez�i:��xF�u�˗����.f'���M
������'���5�g�2
��+�U!��bm�T5+S^'�+�.�v���?��	�%�ݾ+�\,�jc_ɤ�������/�jM��ZUwGS(U�|��?'���ǹ_�]�D
r����{	��"��v<���?Cv]�\����҉�%�O��=�z�Z���{2� �t�37���ǒ6M�����l:���M� X[.�"�A��<=��$R��9|%U�h��d��)��UFA5�n�j2#�q�O�����~"	1N���y��vx�5��Uұn�gh�6~��6*B:��Ք�Q��V&o���/-��It֧w�k2�pi�Z�敉��5[�_5������&�s7^>�����z� �Q$(�E�q����%��S��E�i�y<7�"��oS�С⛼�����������]��{w���OwkU}��E���k$��&-�h#�~���⽩�ÿ�>���z�d����c;�vq?�&��s����5F��ꆐ��k�����J=zᇳ��t^j�ts���)l���r���i\C�ސ��ܗ��/䴅{�KX���,��ڼ�6RM�s3
�/Es���R�1�@tC�WYI܎�Z��P0����W*���ʭ��Z_�G�:t7zպذoUM�.ת��p525�M�Z�뻁&q��)���ɪiO�}������ZO?�G��L�A����?��0�e�?kr�Ԟ��'L�H�,�S��
 �gHG$�-�;����o��_+�h�{�{G����|-~���6R>dv;�-��8eZ�<_'�8�Gc��P��w7 -����;����~2���P�5�"��o��c���J�O�,]��U>;��[�8 (���s�2j���t;ܐ�%�2��ӧ� -�0/�-�^'#��ϥ]h��t%+�|ؐ���S_�T1�u>��]��q�F�W���G"����c7��N[pX�ۯh�(K�(ɯ�0����Ά��GD��u������>� �g�zP~��z,��â�c1S8��~i|w�SJ�����-�B%^M����L�G�Ľ��i�W���s�%��X�?s�	[�4��j&N����u*�vj,ܹe�@��<��qi�2��^|H`�X��gll28��_��1�$�PjJ&Dr<��G	M�eν`�6n�$~!F�̻��2"�(�w@��[7�}7�-�o��8hg��2�Q?:pl	vh\!x�Җ���6��}���QF���p���0�>v�k~G͑o�r&����}eve	n4�!��S8�����?��[{v �`H�E�D�4z��ދ?�i�k������c��ht�f���\��L�S7ƿ����q�[�Xiؕ}���zhq�o~h�H,;W�ML�f�ѯ�E�ʉg�/9,��ؓ��6
���]�]�6#�#!�M����࢈�%���ݸ��� �+-��Ӝ6B˽��f`�6@�&�f}�� ��ﯕ���;���6׶�AE��9�@�w���3D<<�����䰀�FF��AA��������i��@44��b��d��� ���\��,���,�$p�U��Uk�����J��T ���5�͞�G��DW�����}�-'�[��
!HR�ն�����tr��;�/3y���q
��fg�GQN�{r�gh|�Q���d�y��'}�7��k�$�i���T�����H�Z�̂�0�����m8�~�F:�̈́A�)����NU⋮S�*Ϥ����*4���o}�¥�;�
Y�'kr[Qq��T�񣺕�:��+OI����m���[H�����>]�L6Ef��3�����1K�Ԛ��e�b���:�����Iv�p��9�9�Dteg��l�R	<�4�
^�ݠ� �[�����y�ڨ��1Y��:|�}: s�<�9�͈�xW
/n�6 ���#,�eM�� �;�� ��jX&�f�D�E=�/��!�U�����8��]	�7B�w똾k��Z�ț,|�7�"�7��#z||�����-B-  ��Th9W�	噾��P:���,��9���?Ǚ)��w�����EL��b7Y�����]L��������H}{a܍]S&�f��}ul��o�Z[�<6�����F)X2�'Q(Lw��Q�M�Iq�B;U6M����C:��-R�0���3`�I�v@ҍ�4U�V�؍�h)�q���qW�mc��r�zK^�WQ��o��L��t�To�Q�w2rr�C[E�;�Y3LB�eQ�ɶOw(�4]x�-�}j�3�B-�ڱ��g�/���+��U�t���{��Vb/��Pa�jkp~�������!i���%��kA��d�D"wBGc��{�d�)a��^x�[�\�g!���s���@<��͖þ��U�EN}�;�R__�@g�>�._J���P{2(w{|nNBl7���&��Lw�t�M�i���ɡK�-�Pz��:p5���q��Q��0;�ݢ�Z�S7�Rvړ5ǒ�S�pk�ھ�II�+�9p5#�g�C�����z)��^z&�W:��r�-'W�%'$�"�BJ����TBB�����G�TTT�<���␦fcck�}��H���~`��/���P��m}6y���4dtd[_>5]�E[��y��C>���ID�w��Q��3��	����C�-R[����\S��Є�+�Å��L&��I�]��X�n��Cg�J3�=����G�h�b��0��S�l+x��~���0� �Ɏ[�	L�dn �Cxs�_���\���c�>�>��e'Չ��ш:��s��e��'۾�L���@4x:������dS�K��@
%D��k�����B��
����[�偖x7]�h���#�#�	�]�K'�S�����Q���)V
TQJ���B��5l���Ɠ(n?>�G����Jϴ���7Q��C#���-R����q۳�x�L~X�Z�<�r�蝑�Ї�t��s��vW�4��s�M_�=� ��W�ʶ�&F�oh�� Ym;�#'���ȫ*���<�:荭�j�As��I��������唿��ӑ��^fQ����9#�<�L*�j]���Q��6�MqX�$"��l"qg$i$�QG�ה�M�+M��d�^��\��4��<J�(�"]i������A���a��Z7I4�]�'+l7��o�N���z��?�4��*���g�.f�������b������}g�˿���.�m���㘵�_�P�����Ⱨa���JrSi�n��A��j�q���EC�jH݊M��I��n�� 5��_
�|Z� B��OC.3'E��c]6�N��?��Y %��ʊ�ﮍ���%�h��_̍u����I�\?]����z�n���Ҫ;'�otM�H+JpuiQ�6�ׂ{��K-�j0��Z-ؤu����,��j�҂��:��y&	��|�d�}�
%KnnyDe��"��Y��y\�B�j�Ɉ:pK&(�HR�Z��n���T�����sr/�/���2�H�h�����@+=B1P-͙���NE����fS�Fǖ1�>z�/�e9��.}!�;�$�@��'�8S�5�XF�UҼ�?�m��}�֮(���p�35�n�� R8)U-~?�^��t{��'��a���f���I�葳�ϼ��j|;�D��4C��65���Wά�6/��� n���h��V=�߈��M����"����jڤ�õ��#�?н0hgV��I���2hjo�Ѥ�5�dI��0��y��KiM�,w77QV�<��E�iL��zI�9���A��5�±�K��!��jϮ���l�9sk{CC�8xp�q�֫��}�D�H9�ާ��j�,3�[���sˍp!���,>�Ą	,�m�f���\�iŴ�Ԩ�ܕ�n���l��tNi6��u�z¸v��< ǫ�PL�z�%|��3V�u?�P���v�k�ܗ�9N�����a�D[ӳν��/i�	�Q^�C�K��(�{k�	�h���E���-��5f�k���r��ə,g�h΅I�9�[u�a�ޫ��$�WF��� 0�ڷ"���u}�)D�����t�xw�h�bc��Q~
e�DDR4cV��Fk¦\�3�v���"PK�uC�Ƕ�c�u�}����5����)ӣw��B}g�b4)Y��W��Yt�����,cK�W�yp���](t���>t�ٶ�MV���r�W�h�^P�~�T<� �W����N2�ML��k��!�x�J����G�����׿��'>Q=�<���h��(���
7�^�7Co�X�F~b��:ڃRs8wzH1K�u�k�K�m��� w����>��ݡ����X��#�䋥k��&?}�c'��2���W��ɿ^���wO`Y1��\��Y��,��֞����˧S��*U�<0(�x�r{�V�|�%-���m7660	,V �KL0�p��^ױ�������1P���;J�a�4[n$-�����C�P.�SB�t�:%Om����9��W�b8�O D�R�����A������ظ�'���ʱ#1�5v�"QD��O؝����(��`��B|�&b=� ��M�-~�"�
X�_Ҫ�z��R�ɖ�v�k�#��P�sT�"����S}Ev�auN���043���s��ϧ��`X��!��?�K�bygƐ�h�+��>0q���*�Q�����Ow�`�UGu)$��	����͖�2A�S1"��RMÍy������r���lQ.�߇�4���������b��<�j>�We{�+��N�xs
��u��i�SY�Y525�J��e6�{V��hp�(<�<�a���eQ�n�s�3H��i�։PD@3Ț�/����9T!�����;��.e)�J��R͈���$'�O��_Y�J9��8C��1Z�(Ɩ�*Ǘh�p��Ѳ�%S��X䣶?ɀ+>��l%�)p?s��%��f�;�0Mg{�K#�/0dM zu�8n���(�h���>.(�6�t� �>�oblu�tw�U-|'Fa,޳�����+SYI�0IH
Q#�veG���a�И���Bڛ;d���ڈ"�7=���̭���(�b)bi�3�쬊ǜ��ړv춄�54H|���9|e҈O����#~�tϬ���rS0<�gY�s��,�Ey2���E���u9����c�u��>ZTM�j��^}F L���
����M�Ok�'PT�+�f�kk��@4��ժ��ZJw�0;Z�_��?x��-Y�8$q�ڟ�Z,��ZRu�W�|����Oe�\�f�>��ȼ�ͦB6��[�X&��@�h���ܺ3�_��x�#Hq۽��v�-&Y��4��5a���B��iM�Y�w�	��p{���x�� p8�e���s��w���Cj�c���F���aT���j��lY�Z�����T���j��-8zH�b��N�j�f�J��>��n����O|�\"�(U����ǭ~uBcGz%n�c6��o��A����h�i�Z=G_���p���yИ[�My�m�g����ݙ{B���G���ȥ-#�!��/��iMONG>5�~}T-�z<�����-�81xx2Q,r�p�b��塄X:m%���t[秧��А�	�Sh.Yp���VD�b_B֐����x���-�`�����*���G�nARR�NQ����ݩ�tw*ݒ��N�wog�����y���s�9��k}b�u�N�݅��U:?�q�<<p��~�@�|oo�]��RX�\~�r��ŗ/_l��4�hx�+�o}���[rˢ��]��8��lb��Wg��ڬ���@�>�Y&�)4o|�z��8M0���y��M��� P͟1���z�њ����0����_胳�2Oa���|�ȗ~���=o�R�5���N#��k����n(�_�7��r�|/����{���,@j�8ݭ�8��]�ݠ�ճ~񩲻���$�]�` "�ׅ�L��):9��b��We�]�?2��*���ړk/aC��*\v9��/Pj7�����>~&��H��31����.��yS� ��������a'>��#�����&��|��P�cyW�^� MO��X�?�����'�{AP�83���z�8����S_#�އ���``���H-�5�d���俿�D�-A8��r"N'�R7bf��9�|w�:���G�441��&λ���K �,""�.��Z��W�X��l �)7W�����_����=�3�*>G�+˄@y��mm�-���짶��u���^"P����Ю�U��%7����`�j�I K��	�!��!�⸢I�&
L��"�~��U����MN�7w��T���S��s��,*)y�A(��A��ro�i�}��{ֈ{��ZJT�M�j�Ɉ"�8��c���7�������^ؖ�%^Lv���@���^�@T�5>&9�L�sVW�2��c"uť����F �0���y��Z��&����Vzb�`q����цb��&��|
�M�`@�!�U�ra�� wg�<z���$q�)'��~�3S�?�H��n��Q2���u�2{�n�����]m�撂�K6���}���Ve�
������͖��u�����j����)���|��^Bq�m�}֤�J����$���-.*)��U����m4�BԦ��C>�:�B����U<JJ�kX����O���Ѱ�t�:^
�}����3�9��4����(riq?�����n��܎��y���8I;�� t*|3����ue�x�-�Q��@hy�k�7�4���yi�۲����T6d@@�ͪ�)wT���2��"@2U5Li�,��|��#@Qdq#: �(�X�*�>YUxh2�|ȼf��EH��r�8��0����4?S��[��=���p/5.�K�}1���v�~O����(彮./6\�s�,'U�?���,ֺ��3ʷ��L&͊�ڲw�b�)T�7i��e�LZO�
������s�� �s����.tjv������'�dˬ��ʯ�D.C�]����<V������B��9�9Ȳ��{�;å|}��4�X��vµ;�f��Bj��
��A�ecs��E�0��״S�2���^>jג�oA&�k�|B��C,▎&�KO��n�Pyƾ�]�<��{���Þ��>����Gv���I�[��\���$�񜣭_���?����)l����R*�]N�]�Хް��&`^��q�h�.�%����a�Y�=��<M'�X�{K;�]	V�la��<=��a��3r�9��@�q�0P̈́{w�mϽ�6�F�ޟ���]���l�W�8�k��Mg=���Eo�8��?9 �d�Lj��qA4"�":9��|�ݤ�r������o]��jY}򔝼�U�s�;���u��x�3C��D�]nlQ�U����J�J;�&$�x��}����F�w���I�������^ ��M����m�� ���o�*�T��+�F�n�N�Z�:x�]%�o��ܶ#v\3}�,�z�A�Q�l�{(̙�	��s����	)u�Q�8�s�ڨ�J'ؖ5�}l�.;����ܠ<�%����v��P�:�y�yA�>mk:��a���$�q�=����U�~[�6ǴB"�o�ce_�$�4m[`x�u-�G������5a��`�Mf�goq�����h&6��A�f�Ps!ޯ�@(Eh���򺦍�]Y�"�B9�aҗ��ĳ�ʀY\��v ��J�7n�a��*��W@�o,-�e�v� Mta�K&lv�RY�/�Z��^�1	�
c"IS�,G�tt9SI ��;y�;�˵%;�n��g��ѩ����>�D�$�t�y(��BKF���9Uw�]N������IL�/��{&����Ɩ{�[��EY���7.�M�g�5d��S���?��]������
���2��N�-��B�����FW0O[R����]H����*��.�c�i�{�J7w�c�,��eY*��q�3H�U�0w�
4k0m�P	wX+����f�}��v�����S��������᷇p?>��^����l5&�E�v���ngץ��n��f�{�z<�X��#e�iʘц�4}.�w���f���\O:S�j�jG���]t��"���+��DiC#j�m�'L$A��C�8������b���V4�IJE����uM
�3A�<��$�D.3���hD⑿f6���7��YG��5���ë��#mmri2HON?[k#<�g-��qA�x���Khն�l�d�v��XG�~�'�3<~�75��{/S/c���9��y��R}��"�,�˽�O_?����C��#���(��J�W�<6Icd�R[�٫!J�Nᄻ�h��7�G�pP����D�����#�O(�!������#�}i���Ѩum�2��e%pG[��W��=�U�l�\ۅ��p��2��������F��G\��w�js���ڥd㿑��,$Q���F�b��\����s�nмY�fe��^Ty,o5��VRޓ}�o�)�1�f,���G���(��U�\@s�w4�5�04z�3>��z]�g�Y֝�ʿ����v�Y><<�I���&<<|:A/CXXX��	I�T�-mmJ.!o�FS��} [��-4Y��o^��C+�|t{(�*U��&sM�;�A5��ͦ���A��룋�����e~s_�c*� ��0�6�EFR����e��qK���YZ����$��J~�� 9H�_u�gھ�A�>0���A�O	]�^�;X�G�[������M4v��WFE^��_##��lccv���J;�p���
��nIU�{�(T�_��1��m��޺{���'W�V��܇��3S|�k���ux(�z'��X䩎��n�g%}[.�;��z�a�U6�?SO��е�皴�M8�C��.I���o��ـT�{&�$��o�Y5�*j\}���|��>����:�h8y �
��":�����%gs8���3�!�����~���R
��f�ff�ܺ紂��#?x�Po[�Ȏa\�M`�#/;ݷ���4�VG�`9D^ʇ���3�\uJD�,��g�&7�O�D���y���lN�������R�`���Xd��Ҟj�k�jJT�^5a3�Np�58��ǝ-*�g��1���+;��gP�
RdK%&_H�����H��_"�����)ۄ�h3�� �±
*�ٱ23331�i��:�Y�B3�����/}�[�-�l:�{��9w�xSh�n8������IáΙ�d�$qJ��0rp�L�xYÕ\1�������^jhUV�L6�cKY����ؠ����\�mVm���4c�k��l�-��\�*2�5b
p�ςZ�,��^�HD���z��h_��錘����I���U�YAܚ��UØ�&w���38)cŴ]���?lJ=Q�Q�$
�k�R�	Mw4MDb"���!o����j�:y ��B�**�b��d�l����Gl�+��7�8x���猷��<�Q^�Y� ��.#��ɿ�����ز�󥧆za��� �Te�CJ�[�r��Ǡ2�`(�1�Ԛ �F�6E�Q�-���.6�6IҦUt
���J̹u���q���
f��U}Oa@�2e��CAJ��0v�O�sC&�ƽ{�� �aȅI�Oš�0Ԋ��K>�^�p`~�5G���=)b�M"%r�=�R������3�owRп}̔H��*���#�3v�ˣ�	yY�S�N%����$�7�L�V��k*�U.�^'ǽⷿ�[������ږϑ �|�˳�Pd����m � J밭t%�|v�R�!$B5B%#`K���YZ_9Y?���^�������{<���v���-�GSW�F��`���=��r)+9=k���j��g	�
&�С�B����"�YӞ���z�A�����5(�K��ժn~���|���>�z2O2+1zRgVǫ5�J��`�[4�l���[�K���\��޸� =��V$!#�b�X�@��������ˀG�ND��O����z���PtMT����c��}�Kp#���,�h~�$�Q�;8|a���R�F��J���5���<��ۛŴ��J�9ayt����ׅ��ʎ����u���U���P�~ 1�a����J�ܩ����2����׀���x)8W��4f���V_����1<��p�^:ڀ��$-���u��f�ћrH��u98�S��Z�Cd4�R�K��o��Ku���i��H�a�����_�.�������� $z�Ԥq=1F䏙�&�[*�#���|/��q����:z�aN_7-<���+�����e_�Y?�_YQ�����E�"�è��t^�\����������F5�卩gg��˲Gڔ߮��3�Zv:�f:�>��ȱ�CV� ���{i�՟ #�힖d�Χ�R���}DE���?�:�~#)q_'5a�HJŹ2��*m��|�j$����V��oN����Z���o~/��kt��(Fݾ��Z'Nj��II4�Lש��Ǥ»À���^<=�����ҿ�E(�d+�X��y��[�y�{RqT'��L"xnxp�tt�&��l:Z��J-��j�[��G ��Ĩ��Sڟ���F�*��L�B��Ҹ� �����������J���W�ǌR��y7�#"G�_��DG��G����8��y{��np6��\��"&�m�Z�zr�8�@n����Xn9w�������Jms��1P��4�e�i0?Zv��]�P���B�7�a�d榪-?M�	m������ai"�" #�#Ee+���޻7��}�p��N�X��v��M�Kf_ճ�!�Mg���G�������݈S�Y�&f�L��uX-w��쭝r��F��r��W$�R�TF^+k��K���%�"�Wg��C��00
�|�����A6��@�4Zi�&}���rp�������%�j���mϳ��^u��[΋���:"ƒ+���:���m��?Շ��'[*Y�;<W�������Ar�NZ[C���ŵK����1zw�(�.�4��]�C����6�.6��{���oJ�;�f8�tM�LCEF��X����:�6���d0,,W���d�ʯ�Ң������~zj����i)|?���!<��U�;C�t\hh(�U�'�V��g�S��n�4��wk�����������U�s�6������[�8,���l��{"P8�f*CF����_w�x&DD�'t��lҫ4�V�$c2M֍���+rG�^ŕJ�B{����l�9.ތA�S�"�w/Y&���v�pb!��k����Ô�����>�]��*�,�N^\p�˴��Υ+�8?.��N��y+��J�z��;ֻ��c�
�C�4n��јݹ�LR��
�6�F�ʅ�aN_3^!�*ژ}T�z44����c����=��>��ȥ%-V��"��a��5����uf�|"L��<~h���
9K��{Z��c���kWW�1�&�+ ��N��}�W�����;�@�8���Ue�����z�FtU�34ū&�����#���j��Dܕ.��b��KA����"�-7��+Ҩ_���&ҙg���j���TN��ګ=�z�U�_5ݍ��s��h�`��{�!��F�b�dـ����m�&��Z5���0�>Zͅd����+l���al�L��&_����꽟Hf�@�iN�r�ʂ�̷��PK�}Z�w�,e�ځ�N�`����Ȳ|>�5���n����(xx��J��^==�O�=5���~�0Ý>l��h��!��VR�/nmk��?���i���iâ|[n ���pk�Ć=�2��QB�o�j\�*��jDK2	�S�2/��˵`��	*�\��B�de�ۀ��B��a.+�$��ot�P��TYOa��vl��t��Ά%���0��z2y�DH��('(/̄t�=J�T�z~�^{�Ѻ�Q��Lyz����N��n|5���+�������8�JۚiC^�s'�,��E|[�{?�
<�a���E*�Li�IW����.q'75v1�hV��K�R��ot��f�쌌ȴd=��r�ADd<$$$M����|��'�OH�"#1DDE�j2�l�FCG'cg�4!����ދ噅����gj��l���_�hUvGQ��y ��[j��am��=�=���uAi_�X�w�LO@��+Ă=\�t�X�SAi��ԭ�9��q�%o�$^�n�j��ƅ�'/M��Ȁ�wR;o�a����8�8���C{�u1�XeK;�P�!p�$Y�2����b,�i�4HՍWm�qI����ǜY� �iͮ;�e^e�_���ty��8�!cc0G�
̘*�v6��P#�T3��f��Ib{?�sЫ��4�ċ�޲��81Jݮ��w�4 j��Y�6���5�=�.?
]�|�
�M����aF�`��K�����~00�yJN�����S���8F���p��I�ܰa_W��)Ԏ����v�]%R��\��������+�[6�p07�$>Y0#Dܚ��Z�Rq�V:��:��^h~��$mNR�[���
�YM'��w��F��s�0���w}��VGg�^¤/�.��tw�<�~t^�����y��6��Bs�H������N�m%��h�:t����ʕӁ�FWsS�u�+��dɬ�8@xYV��5}�-$v��|cexy�8��;��&�	@_1_�۽�?�s:�����w������q���������9߶\�.\W�VK5�[�R}d���¡d�'�E^�.O��0U���)�=�w��ʹ�L� \.""���t���t�ǈ�vGOO�sRkK�Ҹ{�M�ׯ�^�&���wُyyy��-�����\�����Ёc
�:��$ �T`h�Ĕ7(�ѷru��>d���/��!�֧��F\"4Z[�ꡱA�!�0���S�qs'_u�,�s^+Q��.�(�W$
�#�#�9��,��۽6L�A��%?o��ȣ�@�e����q��&LH���`�.�僪BF���r0����@U�kĵ�����|�wM����xE���	W	k���[��+ױ}��d-��F�5����3�܁�E�'��_;A�4r`��!]���M�qY���Y�C�=�US6Y9�h�e��ec`��x��?���2�<fe�/���uؐ/��t�8.�����64*J�q�!�G�J����WLK+�M�k�����" �ix�V�~D%�����<&��38�>S��Ap��fo}C1s�
���C�p���+-֫6m;��~�:����}^bpC��mU��F�,f<�|�(
��kb1y�T�T������묷�݉ۖ?C�/2`�D��Q��^q�%��D*�C��#wx�7��K�K���$F�޻&��K�,�>�	@Ç"(��G҃� �Ν;��H�,e��X@�~�7Wnh���ፆ��u��k���������Ҽ�̴L��}-��H�;]}��a�<��}@���:Ar�s s�O&�"�^�Rro�e75���FDܯ�m���A�m�l�b����z��Qr;�(¡�?������C��V����1�di:A��B��N�_��]�O�o�'۩^�3g�����Oc:1<2�ZZ������Kګ{I&�fPU���y]����S9�r���8���! Rf�GZ!��.S[�~���E���x��q���[ XZ�.,	w�����P)x@�SX�W��
�13Ā�<����KUZ&7����5.�]�[G;�1Gp�:ty��Fm��A_1-���aҌ�Y&G��8�ck�a���+��4��z
���O&�_�8n�J2�;ߋ,��#��}�W���h�	������Q�!naq��JǕ[G�֗b�+?��>r�8�n%<h�!����$����*�ߟA5�FX�Vxx8 I_���նJ����(��̞�o�����]*�f��h�v�]*wL��Ȧ�Ad���x��ŕ^��}x���� ?R�`��ۂ7����w75�:�9m_�.��4D��h��279��!�9�r��Y�}m6�60�	�T�dA�b��dC�(oT�FJc�=�֬���R����̪a�~���|M�a�` �˷O�uK�+��^4ᔞ�L����ƅ��,��q	~�C+O.1.N߫���]LE%Q/5��Ay�IA����%�� BQLA!VOO�<��i�ֹ��*,�� �#�G�oZ�k#������={��7�Z��H��;�I�'��j���7[2�G�����[��)���������;�(Vm�
�`|�qbz�01l��=w�#��.���O���?p9*L��\��I�r.�ks�܍O5[dH����y$=��, X��U��m��i��z��ہ̣�+3�D�YUO��>�c1ҳ}�����վ&�lx��D|^\\\�E��
wh�YH3n��g0�s������;� �/�O� IM ��-����o&�� SL��:a�Q�p�)=JAz��a�	���tEG,�4��.�7%�#��a��g����S��8���l�,� �2\xx.�9!��:���`��߬#+�XZ���P�J��M�ˊ�.��A������
���e89�~49���RY�^(��ѷ�����Օ�]ʞ`����/����WK�zΓ�Z=K������ʘhXXFM��̊��Ԕ��H�'+��j�MP0��H�,bx~��˹ �d�|h����*)����l'&�*)@�	��}�3�����,>�m�졊�tF����j?����n�>"�yUjY�����Dc����Y�7Y�YJdϖ� ��pH���PI�����K��H݊'h�Wꦬ�}�w��12K�:t��k����:Ld��︕V���	C���I�t��Ә�v&�d���{R�+}�������i�D��X�A�xV ������b��$����X�f�1�sp�a���J���f�v����Mg���ɜm&�l�+�O))��;q�À@%ڣǹ]����F�`�I]��H#I�����k⣘E�������B�+����謆�فoa`B�*�IY/��r'�Y	k�h�ӓn��g�j�h=�_�y��CEȨ��S��,�A��ۼ�V�奏�����+"��;�8�>����ݝ�@�(��3:ŸK�ɥ{>t�_�wmpw��ֵ�I����Ɇ	����y���J\�g~�\����+EA����i'��n�G��t���@/e��Wo�j^��������E�����԰�Ild).�ف8�|�̌�0e8��ذ]��ӳ='_U�������n��Y@n�wmU��^*�����	V@��粧!W�r�W�qk���V.��q����5*8k$<`<���� j{5⳯T���T��b	����&��D����'!�J�
H>�{t�!�Ï��`�"e����67<,�tv�Rn�K���$f�Ea�j�����r]��`���y�����|,���;�W*�*�֡U)�/Tu}m�h3���H˵&���� ��pn-<>�����G{�):6��0ٳg�>��(<s7����ƕ�Ϭ7n��T䊋���H���~��,oUq>	"(�6|�S����7�I�nΪKܕT2'S��Id��ջ�K̛��7�e�o���^�7(f�i�],�0����k�Qq�����0�/�/��==Y��ZmH���'��W� �|FGk?0������撲�- �)��U�:s�zy���%^�vx��Qh,�)>+w�s��h�0��{�	�5���͛76콝�a����_P���$5h !.f�
8�қ@��y
�}�~�QR��6["D9�ۋ%�~>q�Y�;�#��`צ��e���F�Œ��s��z�e��]�2BRc���|�|��(��v^�� ���K��������j�U�ü���8� ܿE�p`��A�S�'G���l���31;�'�wr�2�8&VM|3���&(����
�8 ci�hhz�����b�eddL>�T[���������z�1���EUH��+�0*��&oOÛ"�9�s�����R�K/1�exR�87����2i2H��!�Q�������bnj�Y)BX2:͜%K�`�9�N��ɒ��@���B�ZӘ�FW&��Q�������?I	awM����H��⑔�b�7��L�-�bպ3�L{��WG"6ڭ4�tm$+P04E��	&<��h��,`C����� ����G"�7���T�+P�~�����b��ܥ$�w�XW��շ�͂vd���y/�1=\9�I�͝e��Hy-�e^�9	��L@�E�H7d8ưY�eT�w]Q�Ǘ����m)��Ԃ�T��1�о�s��_p��:�]<Z8�C�7��^���)ٸ������˘m<w��B�Y�ݽ ���e�rX�'�����p�^�Ǐ���3RQuÇ4�zyyMI�N� %|$��9O���̲Zl���5��H�l^s՜eó���n5<,x�
Վ2��U���)�h�=�(���%��s���:���ϑ�Y9���,���nm����OIi�"*9�X�Z��DM		K�uM��f1w�ܻv�����usſqq�؟1��VfY� �_�����A�	����v���k�VK��_���~��cJs*���U2 �`���"� T�/����Ad2�x'B�:\[>�����
 �e ��.v}��;�[S�U�-L�^��' �3[
�W��լ���ۊ�!>�z�������:kU�kCA�+�O��h���i���v���^-�Ȳ����i�]�v74����MKN+��5#7��R<]�.ZQp��8���j��W���I��'�b��'?�r��:{�z��m\�w�#����bUq�����>������a:���1� X>>��/s-�/�p���p �<��I�`zŮ(��c��V�n�8��k��7?��caD$��>�>|�teA +=<�&��fV�]�0�h�k�kl���)F��c�����a�ZA[���_��d���\�-Vך�j+x�<�� �����i"�c(eg��fƷ�Lc��fo�M��rwm�b���V��)�`m��@��ậ�^��j�a�'{x@+��84֣�������/$$��E>>���V\k�II�,�l��p���O��e)���Ƴ`�O�:Y��ö*4I���,�.<*xT�u�eY�q˦�F
mm�x���dR�S���N+��n�B���E{�!XK��]dW5>O>ģ�Cj�X�W�9@�ơ�4���N�ƾ@-6�#���;�4�`�:�M�}x�?�c�a�nW9�l:����*�lE�{r�UïX#5�5M��Ô���S�H�M�,�/X��Z~Lp��w\]]�>|x��[���{�s�)RDR�e'��R�V��=s�9������#����CX�n??�]�H��'k��_-a:2�2z2�lO'ڷj���3�u��u3B�|�A��0�ן�_�.���^7����ƚ�Etn>s��Y���c+���۹$	Hv�����'�?��p?�Ӭ�&�$�Upl��d��ӧ��7]�����}�� �^�tW2��(��BtM1����X"h�M#�{�9�m�}���`��[�8�w�-3ԣ|�򧓾 v��1o8D��V�#\���n'���pF̦]�1ƞ�B���Q�5��f�_��Jc� Z`�P���Ѱ�ɟ?ޖYY.ɯs��䒙*��^��1(
�n��y�S��{,���9X�Z94F���g>4f-+��d��G��FE�6�zJ+_�h��!3�^�=�E�I�ܴz�q�Rø�Vi���;������h4TTu#$�	�o,TTb �|ǹ�G �E� �|؏��!|$��y�.�[Ǯ��!\:�ɇظP.�+���d�vI�vv߅D�G>��1�Ɩ�[��IU|W��,��)�|Ê�x�{9��e��`ЕC�O�Y��_��,�c�]:Ԫlg�7*��\����⩕w�ۡ�!�x`�g���ҳ���2��eh��;.v��n?zw5�=�C��������i5@�-�����ת�Þ�_��lJ"��j+���㖼�I��~��nY���2��Ar�������lg��yOM'?����g��V��@�g���hhh�<qKKZO�w7Y�0`E�S`�Q��n/���oж0�4�VjMS��[��M1=S	~J��s*	�m=��S��N_}/��;�Ե�ںNo�$2{3�����w�����O�l�{��}�?��� �l�6� m�F���ö����������
^�$�<
�[>"���玐	�H	�z��yl���-�B�+�X�9�]�ջ� ,���mS�V�q
Q<��/!x�ش]�$�
���#������������)��TO��XZZ�Id�탏2	x6"�⑈ش�\8��[��Y �{t�bN�v�X�qY�T�(���Ĵc���4W�Ե\���-�?x���մE�}����1B��'�0_X0��G?�7��RS�SR�<���U��k��o�La>��HQ`ះj1�0F��Xn�>��{:�1�x��ݪ=h�=���8H�m��lN�a��Z�7�\ՙ����B�+M�l*W�{jv���w��N�_^0���B���ۯ��ڝՒ�������-����QЧO����B�шJ��*�ٙ?ug������jb�d�$�3	��\���Fu����Av�a�p>�JA��OvmS��M��["M%�rs�TK�ˋ�V��"Fʇ����H�-�88��Ϯ+=M��eDб�W����d�+������5�m���q����jI�����KI!����n�mkk�������Óٍh�4GY��Kϙ�O�׫7�<��_����:L�����1oi��ym&=�_�"3���Bm�V\}o�u�*��*;{p��g=c�^�x���a���誋��Z�Q���PHB�y�.K�����5� HdTTF_�E��H����z-BX��K��J���0���un�}H!� *
FDp8�_����UM��f�m���^��(V�q%s2\+ժ�(���E�DY"_����')]_����I!�b,:�����q�i�y�9m�_������p
�.�3u�f�y�?���$Ԭ%**�!�"�DUc`b"����=2�w����ªe*w����OBn�BB]�Z�������Xա�����e�����[�"�sC���PG���Ɛi�u#T�!N��B�7�N'�#3��bJ1����!�������}�_�ؖ�F��+�����8Yb�8e׸w%�b��mO�Rj�dk8��UZ֋mB��Ѯ5���<�G��.��(hh���5^�\:����r>'��$g���'��6Y�Cb�H��@�}uw�3����	_�bO��Ե �@��0S�t8�b8:�3{�;�O7kZ�yЧ�*jr�@^��MG�����X_�h>�۴E�p�se�7y���^�����h �U��[����д(+�̘>���>��v�U�j�U�fZp<�Ĥ�>��3Ev���Dw�Bz'������b�Ǫ��'i,&.�+z�����_M�o0�B�!C���W�ñ{��{�ƍ(���7a�	!a 4�#�|��+p�l��6�r&/4��f�N�z�|n��`�6L�˱�)/�?�C�b<`=I�|r�4Z���R�#���~f����r��5�\��q��n���Y� ����)�-@�2�.�fN_�~%}�F&���{�i�%�����GzU��o����3�p�5	�-�+�Nk�&���WY��J'.�5���R�)p6����+�{#I��I
�?q�޿s{5��/�"�3���0R����x-�b���UN˪&��փ�|���Y9^D�$1޸�ތ��e�}fb@�VoC*�3Vd1���E-�r�^��ja����]�ğp~�5O���P"�S�@N�l�&�y�;�\�.�5%��NN�n���4��_��)mR���I�媱���`/�d�w��ٯ��꫓&��ɔK�c�t��/`}*�_ou+V"`�\��N:���#Xi�j�j��'���f��b/`[�	TVjt�3H�_X>Q���!~�i!.��L�o|����!�/0;dblr5ew���/ ��T��m�%T��m@N�HԹ�j�Rn����;<)�RK��t`������?+��;��J�:y��9�<�Rc!<�d���f��'C&C�+��f(��U�5���r^�M��{ʹ�V՗`��&����V�l�V�[Y��M��9��	�	>ROw�(��wi;�H����U��k�ۂ]x�!gB�4n�D��pT�wE�E���G��(�k	�e�B��Z$�aKU�z��e޻!q����37��;r��*�֔�7 �%9H��T&p�{�i�	M�wF�G��ߠM��r�m�(�7qyӆt�{��EZI������O�#�C&�Ŋ!����J�j$g/�ug�=��|�`����R���4���=c�m0i3_���I����G�a�Z{?��y
<-"&��^��]��`�Ia]e�=� ��fW�3f�<)%�Z�C�V����aB���2ߟ��M+_9��Q)��fN�m�T�?A��b׻��(��~�E��WEb�l��ޕ��Ҥ��d��c
f��C�m�?�:5=]����0��ȼ�>�0�{�J6�[4v㪡�̮��W�)5u���{�D/C�T��]*+L�4c��?%�1����?��cա������joM��8����G���"��,ԙ��7�-ƜW��E��e�$�j�B���J3�щ*�d�����7ҧϓ5O p�|��t�˥��f�T�)�W��6��*��9�2���ܨ�o=	�8!|9E�Ϣ�r��gh*�+����N˷��p
Uwʢ� �դ}Qα�O/��D�(����{�!�v�W1��'n���  �9oN�q[8������hb!u��j{��\DJ�_۸{T)f����2_4�{�1V.���ֽ;���xd�%�ݰ�C���Ar��O�ה�!w�=������}YGl
�K�r�f����m���\Ok�`�h��x������vN]]��C%��@2;�ٿ{mB>��0-c�˚@ ����|�>��E�ׅ��`HJ�M���W��x^Й��T����8n0'u.RJ������( ~ �~C��Һ-��h:�u`�8	���o!�x�eJ��-�R-��eCUZ��eR�J��͓��0%b�z���X���$�m؟�,@��D����k��Z9׹�B���XLt�#�k�Vc�V�S�[���CbGY
�k�6J�?W��z4u�T6�(�H�C��o��=88��{�}vc�ɣ��Ú�?�=���BGy��[럅:�	*;*+��ZV_V�|\��p+�	�q��X����ic�՘�gn 4�P
��:��L����G���@�1�ɖ���E��(�S>�U���m�~�nRA��e�__Y�x����d�k@�.���������U���ߎs,��eb���]�gbޖ��>r}�:�8=a;��{��p�2�L�n��q�@�e������=����g������� *�<��uD�U{��Cɛ-IR�BD4u<��-�������5�Ĵ�N��ij]Z$�B)�fq�5]6f[��O��~Ӄ��	#�Pmml���U֒8�a1�l�U��K��*��@��MLL*i��׶���F��`I8��[g�[w��KV��#��2q���\�n[Z|��E�_y��s��w�+���#��֧�#���W�6�Ҡ�tO�iXʪ��b}���x*�e�J�tŽ[��ne���b���8��������LGfO��r�ͬ�I�eG�:��nK��&-��-F���I#�(�TÅ��Ѹ�@��.=e��Q�Pʧ�,{1�g�-;w�1�������k)�E�[�w�=7S5�-ev�г���;�P���@�r�Sq8͸�@���O���e!�LxԪLi��
�[���HC���_�����9��!�odh �[�ꟽ�9	��uݭ<>�k���Ac�`�ϗ}'��=�ۮ?��9�v�kd�"\:��q��A +h.]�5�t���b��Yҩ�fN��&㙌e�l˲T���[��N��R?	�'�=����2����G�K�q��[����-���BF�6�,�\��
3u�4Igٌ���ie��&-�Va�ϼ�j�]�onm��Z�!j�8�N�&k��ܜ��Ⱦ�e��{�p�&�p�����)H�a!�Dk,n�����igKJ�l��(�f��*��v:�V�5���8�Ԥd�pm]��NG�f7��{��5K�� P�����D����a�����T��.L�i�cVi��$���,x/,x����߄��D�BIvLF�(17�"�,����͉����ɍ;ԟHt8I�PQ5
�*�$�q�"�6�/ϥ�Z@�n��ͨ�u��fXJ�L�S�I�ů��zΝ�9^�A`���F�ش��F�$�ה�����~`����JV�&D�2p�w)TM�m�f�r��X�|��I+\J5	�����7�box�\��ޠ"����]Н0V� ���Zrgh^�UJ�����P�c�*{�$�"�⤿�*�9e�6��bY�`��j �|o/$�����[!��8U�&T-�8ֈB�x|H-�rtF�UL�C��VKJj�Ɂ7}�Y�^��z��q߂�Cz�u�RBʩ��馋�H]lN��]�y�=h��x��������;�?�PX�R��Rv˰B��$�d{
��X�f�	`T�_]UL����d����ts19b�/�e*:ک�`�d1�^?�:�t�m���!������ң����v�+�����v��VF���5~Y`A�A�#޹h��W�VE�ٛ<�����BQ��>�h���>�����r��X�l��~"����;A��Ҫ��
h̬��k�m���k�)����fK��G��Ī�N�̡�]�Ն'�n)�C��Y:}��m�s���#�$)�����s����y����u�¢ ��aH-��ٌ��n�L�O���l�� ��|������*hb�dgq��o��a�]�q���v� �P���Y�s�6~���'t�6�ki�?��:����U$��P��n$������
J
H���t�Ơ;�C��c÷�G�s���>�~����s�5���c�9���7��ݍ�a鷼�3fbF9r%��7ͥ��Z�Bq�+R(�	��+uYV�ţ��]��L����Ⱦ��oΔt�'/,%���E�)v�ojn�H��U�1�C�pC�&�F��R�l���$4�L{7�6ħ����b��.��ȋ�PsW��v!0e�_#��]�Έ��0�J����<�Q4����A�$)U���j�#f����w��R�畴}��ktE��bl.�b�y=���gʏ����Հ>�ȿL�?*��&��s��iW46�1<��5�˲�֟��f������m]k1)�n�)_0]H�\����̎Wrٔ���Ï�� L��ا"�7㽵1���'��g5�1b���g�P!d�����j�#��b4eAt�¥��-7��KC���@(g��Q�p��3~��ɞ��� �_1T@R,��tv�a�k��e);��u�=�f��X�$M"���8�{Nv�� 2�ʨ��
??�Z b��V�^u\l�{����Z���{x	3.����䕃�jꏔ�/����{�^g���\��ͫQ2�C[�p�)�&w��iO�ЂY�{.���I�?���]ە��q={`ji�6�J�{R���d��T��������U�qL戨ӱ�tTǗE6Ġ/������ώ4��-vC�6M7z���̣���Ѕ��o�K=-�h9X�iE�s1z��E]�����a�ۼD{�W�Q%iz���# dӼ3���Gܹ�9�&]����	y;Vw����M���y� �(�f�tGg�t�WS~��Z� +O�F'.�IS�%�]�X	*�|}�%��U�UXD��Dv]o��}�zn�"�N�7�K|$�7{Zo�fњ����jEk����	���.�N�����Y�rם{{GH;�b�N��0ƕ��N�~۱�s�]��"A5��O#(�1&����+����\Xy/dH||����Ϋ�T�į���'��u�eo��.�7���|nT�w����ff�^����C�v�2\}5�I��WZz����(]Hl�!;��E�b�>5���f���a����9�;v�G+O��;t�ʽ���/pD qZ�`2v��{�r��}hĠ��+�x����5�����fqeś̞�l�/����J���18L�U;�7B�4�\� ��n�,����ﮒ""�}W\�3,Ŏ.�Z��w#����-��ٹ�6:aL�2  u^�}����2@�WBy�CïHsR�q��n�B��P��v�������`~�Ar��0�Dk�:o��[�s�����z�./�����3����������q���w�uįL۔W=r�[��N�pZ�.�-AǍ�@.U�P���=��H�M=H����2�ˎ#㣕ykrD%_�[�\B��vw�܌�l=�V���^Nq�fL�3��i�<�C��::.��&j��N9礵����i��O�̷7'Z��<�-v��H��l���R��=y�!�㫎C)wLu��
�g_~h��ƠA��#B��2��K���"�:����*=�P�v#�
����.��"y.�@� �~ވ|�z�,Q���ʚp�u�j�`Uj�<���<��ޙQT<��B��yF����j���ER9`�	�f�ۍ�7�
��V�Ze.�k�E9�w�[*>N2�**e�x3/S�.Q~��UY��M���KKgx�"���K"�z}6r�*��+5�zZT��R|%�nTr��Y�T�?@�(�_W�2�44''cJp]Zi0)j?�P��@�e3;�>��o뺎��;y *My��3�Dd�	Y�����An����{.� ss]�\�^�z.�����F�A|g���iwe�־���H�W�2��=�:�]��hm��&z[�`9�b�����Ⱋ���\L,z��J����EO�@�(�Ӣ��&��qo疅dkf�@�%X�ډ�j��I�oNHI=��i����m��ͪ�E�v���c7�8��z���ǻu���'���-�x�pv�n�qaIX�]Z�1o"����_e������IJS.�{^p��3=��7�֋%�]�֏��R$2�_EJ���"��+�llt��!b�j���fZ�&����uN�h���zXu����5B��#�'55{�C���[�s�����~'�І&�����G�\����A�})�=��"c=����K�
��.���C��$^�m�O�N~ؘF��X_�h��sc��g��Iã8vWڢ��%|�sۣ�~���o�E�����.���[�jt�d|1�yN�_z�|��w➊�R��r�;�0��׾+~���9�lli�ú�h7V�w5C��3��/<>�^�m��K <�U4����zR�*[���K�q��2�r�)��^Y�q���2�o��B{��y#=ڒ��=M��-���K�I�t���^����?'=�fـirR��-���� �����',--��ΞPJ�dxa�,�����)v�ZD\��B�V��L����Q"C�"L���z߿ƙ5y�M��ut-6�3�hK쟻��bj��e�^��:��ť��kW�Lg  ��i��%\쯜�%K��J�<��<v�ªx�S2��#�7y�_?'���?<::z�c�6T��А#��[2\ZL˱:�˘� �sV�����uٮ���f��t�\踰�5�ڰъ��]��e]6WZ�K��)q�p�O~�y�a�VI;[G���W\A�[s���~���Ą:B5��{bFƆ���{�m�)�����_����.nLz:�5� �j]K�hl\��ZE,o<�g�x($N�������Q��Mme�7����ߥ����M�rbh�5p66O����t,S���
��R>�����F]�C#�"��a(�����K��׵�F����zU�e- y~f��1��P���D��{���H�իW�4�C�Q�o�ُ����C����~w)��yX*ƿ���4aNB M������Z�E�޳j(%#��N�2+����Do��-l�wD��p����>g+d+�YLL��(������'ś]*?�9�G��ހ�M���9^���GP�g���֦ވKJ��A�VW'Y�UE�$B�T"�\~2؁��Ml��G�oZ�?��}�ڎ�R9gf�Ar���V��N7&��}��Uq J�G��j�EF�n�9�owǵRS��%����<�k�����Zf����E�o/$ؑI�ʽ�p �4�J�T!����8�M{ c�ڻ<q���hL;�����i�d���h��Fw��7/[W�|��n.�!��W*�E�E�?���i�5X���.y��7U���h-đ��)��\�wt�Եj�n�0�^�&���R��c/�`MƜ�)i�B9yy����f/Vԕ�'1a.�y���YG"e�x�@� �o�Xe� =�}��u��g�:~���b;Q�Xd9��%��]��2�8�����	�R������pK�e�Td���£li�Vޣ������GT7E��Y�qvv��v��`!0�=��݁.QhOqKk/-i�V�+6�`=���.���Ɓ��^�3p���vc��-M�ӎ�����&ۂ�����͇3�H|�����Ǐ�1�;w��f�d؈m�Dԏ� 1w��_߁�������ˑ�Y����5��=Xx��W������!�[�T�l�o��zw��I�Dϒ����3���|���d0Ŗ�8�?�LS��jb�ZS���@[�ڭ���K�z��Ja� ja(*��)��3�
�ɲoN�wNR�m��b�bCX�g���$f)����զ��~b�����E�a \����0�G%�<P2�(G��]�J"=� �?�h�����b�*�ij��͖^B@H�Yʁb�F���g�^��P���f���h5���Py"c�����t�%F]���5�9)�&��Ldy,/-usE�u �?�j:`�1ш񍯉�a��o�*�mv�G�,n�ul[��(m���/ˍk�N���W�خlv��nz�O��I��i�f!��{n�ro �	}�]�
b�5I%����.�\ވ�M}7->�!���h`�m�k���te��m�dP�������lP�c��� �
�=	t���[���R���T;���M�@� ��A�t����/ڳ����z��b23o޿_N���� ��UA�������6DY��:����F4Î���n%�mX�K�iiA��>$�|~�kU|�h���V0M?�J��Q���i3�dI۾}�kY�Z���{-�B��Ϭ+v�A7�`d�A~��:Ղ�0����׆�@`�x�G�S���Y���I�SR��|�������J�s�'�}�|����@M!�GDh�L�XQQ���|3����T�tn�L���7zdat7-�J��$P��^b&ݻW3�%��.�$����ܘ�{P���|��͕���^ە�VND���%� ��3�_�ϟ�V�`}%h���񶲲2 �;���S�K\h���О�<&��i)��^&ώ��iY��P6[k:��y��|3C�����N���C��놶���Ö�-O#��y\7LSF�t����*��w�C��'s���k���ӝ6��}V\�Y,�zzD	d�La�f�_���t�DG�W�����`�����D�)�4�s�H5S�isX�O�x�V!ͩ�x����,�����jgqKs���� o�@/5�mS�]\0���Q{=�����t-R��\�ж���@�0 !���W�� ���6�	9�7&8�m:zt�	����?XHer�o�0����Ė�����CQ�s/x]���,��k��W�nx+K�V�u�Q���/�	/.(_X��8,D�	`�s�<�.R�x*�X���˨=�(�� F�?"'!�����Y�������W���/��4_��K@��}M�R��-�M$��ea:�ڵ�NAK��]0lh�u�p��zA�ѹaecR���>�Z����yu��Ą��݇ �M㈳�z����NZH&���'ERr����#RR*�3�q�ۣL�1t�#��&.�j蟟�0����h&>'��5���4f���β9B5�������y��XAAc��z$��Mf��#Rtr2u>"Ĭ!k����G�ך�.Q�=otc�RS�7Tf�%��t��>�0e~vq6�#�_��n��YZ�^�
y�)�E|m3��ePY}f7Q�Y�#�v�H��mng+2c�C�����~چh�޵c-��m�4�G�`L���%��3��������EH��9[ UZV��8[�(�7cЃ��Lw{ ۗZH�[a�)���!az�ڨ|Z���XPB%۴qkܜ�y�˶����
߁�M�uq�m�X�`���=G�-7"�����_g���ST��>(f�fR��xXڻ%SP�����Ԅ����J���z{D����jEذ��Q��ٳZw�� �!#'�hpM����bLF�3߳^��� ��hٴ�/�y6=�
��T�߫Jx���s�x����&{&4�(�\�J�k�����S6WSS۱��T�5H�H�&�[o&(���ʾ@3�C�S���hn"n�YL8��C�X�--�))��eO����T/�"��k2�P�yuT�pX|ڄ�R� ��x���6�g�gy^�B���;���M[�3�V⪗��.��$0DЕk'WV��^t4͵U.\�S~�������@.�9#�3L1�S���g����?Cǻh)[v"
����,�0�vEʻ�8ׯ_w���h�P�Nîf�@�˄�z��WB���q^��('S�9ݶfp���edhc�h�7<�U��굼�4�=�/p��h]�k]��]��74�^"B>,'�������-�8����&'{�����ˈ=�Yt�X�$%%�+,䢦��NZ����b�eg�GD,�	j�< C�P�"x����<��n���Q��|~n���)�D�1��� ЭR
V��!�r��..�����9�q�1�a���c��h� �B�w�rs�V]�sF���l�-|R�_���b�� N=�u˧���U���Y��')�#�@������v�#3Ļ�^���[��0�-vT�K`z��vC��7�b�Q|9�]
�$���{Ϲ�Y��e*5f�R�®�v�-�g$A�  $�d�q��eP{s�C�F����w�����TTT�"/� �u*�9c5�����7ݓ[O+����n�k@9Ș)f��i7���I�r���<�e�F�[����]߻	V�8�mWn�8�z&���w����Ƕ_�{\e��C&�1h�HE��B��@�|�FXHH$G����5�gϞI������m� �и;w��W�g��E���6����Q��2�iK�����0���y��u�pw͏��\��;M����G.j.D���n�rAe"���9�ڞ�J�������"���C��� �fae�#$���1�۶G�??C���a�M0F(` Q�Y�� 0��+�Kjkka��΢zU�T��q��|���gX۝/�ۯ{�����0�3O��FUlW�]S�et�Jg�^����"�yaʁ�}:��C�=.d`�gg��a��MpQ��zUʼqz�����Cf�\�8������3�!�S[[���o@8���fz�����������
g���*�Zl~�ݓ���Oo"�`�XԱV~���P���].Z�Km�����)#�v��u���/��m�y�K�9b~;�;��N3�Q���q�zQ����A7Z��]���Gd�+���$��~���g��9��Y)� ����|^3�CD�L�,��#R����Ҕ+��o$�A,\�g��%�����X:�N�Oe��"-�P�Y�H��=*���
�^��;��%�ƙ�wa�Oqf���!U
ͫl����{�p�� /��Kwş�_��K]�'��zt1�&|t�MD���ךz{��t뽺���D)g�TG>�xUv
瞛55�C@��<�AH<]h�CP� ��K�9�����s�C�r��	弍���z�:����D$/�=XYj��>\1n:�Y_�!����f2*��ĉn'����_A(//xZJ����<�!rOLP�S;c:��0>������q���	�u  ��H�?J�7�'f���)�8$,.M]��a�C���X��ִv�GE� ~�%@B��A�f�a�n���d�ғރ��	����յ�s��F;e)��k���wL+�r��Ś+�3����k��M������������/����������L#UT��j�Ol�3�Ą	�,﯆ }9��S�c^A���$zG{g�It�2	���}W�M��6���"�_���V�+�<����c�fp�>��h�Z�j��W�^ݶ�^��Q�|����LB;��~
\�~B��rk��З՞7�on���B���o6)�����]��x���?��?�0-�5�z�Gt�)�P���?L>�]�M��J���s��hF W:�P^!��v̢I*4�Ip��z�4O��[+b�C<�ν>'w`��7��zm��23kg���hظ��n�+�>�Hr�MD�r�
"�Jꓽ��Դ����A�;Xh����E}�z�)��-�a�:X����b�C��R+C�٤|�1��+������"]���P�����N^���=1)�3L_�u��Eb���B�%=?o��\ �U�4�|<d�貰�����S��^JE���k�[	�t�m����*\�§�q���%�����;��_������$8884_@�^�L����x��@��p2U��Rͼ�=x]�E���r�G;'�J�h���3�$����R�Ǳ�81�`.W|f/�MC;,�@ |׳u/��@���3��3(@"c�q׸�O|��,�-)��:�i��?♹�9�H�����Z;�\F6:���<�&���=���\,{ɡ���yH� �A@X8�`!p�ڎMvN^JX��!m�EYo�%J��1�<"���l�Ml
{^��t�.>4�*I@;<4jJ�S��!�����z&s��uO�����W��}E@BB�RS+�y*`v�\hn�9-a��]к�L�h�8�~=��C��鸐��v}SSu��ěxD�UU�T�F�L��2�o�(Y�NAN��,�j׎�Ru�PQ_L�Ee���P�2"���ޜ�<�\꣯q���������z f�����������U�2�9ѻ�����64bЀ1�M]�̷��\�cDH��6� �(X�;�ތ�Ok�F���B�  �RSşA?�>�}�j���� �jxx���j��
hjj�
����M4�j}~1�i9���M+�6��ISH��5j|R�j�_��i�������mNN���u�а��o��z�:�7���}�8ozy{� �^C ��r��4����$­�&z�|�di+C�۬ࡍ��2���> !Ԙ���?Z=�G��1=s���N>8H�)?��*{ߤL̇T8[eeq�] ۊ��ǖT�,��n��A#�4�^� Fd���z��� *���:/Ұ�%.�yu���߇�K:>���������vjze�M�K�/��#��H���|����J����
��@�MGh��� 檋WZD9���hi}233e6jAS�
 hM]��.CR�l� �k����������>W��(ݵ /��I�RH�J���ꃅc$���Hx����%@���ɟ/�~�sNf�CZS[�}gCTGGg�z��l)�^~_��8�m���{��i 
`�f����_��d�!ಚ Bs��Ȫ��QSS���H��1��HM����!���j��9a�j��� 	xZ�Ă��ʻ�ӃK?fxի�D/^o�І���q��M%��m.��;��w�����F5�q@ݮ���o�XPl�s���NZY�旡��$|���ɣ�
�&��D~��UUKnb `���[%���ɶ]�9P�����=��9��Z�'��?ۻ/����&�<d�@u�����!���dUHoIc>�2t{�Ɏ^�-Hzy6)��[��ͫ�e��d>|�z~F��94r��hdh��f39�%E�͗�c5f�r���,G��ku��a�_��]	�_�/��aֆ��a:e0D�mzzZ����x����o���h*��`�C�*�#4X1��y�g�M�?���( .)|;��?F�!�M��2��orb���b�]8��/�/hQR����F3 �/te	��b�A
n{O4���ܠ޾FJE.k�
^ss
"�������.#���/���rqR'Jy��'Jy��'J��R��"ػ�rߍ����E;���{���1::��{�V��4�<��7����l�'���K����Τ�����@A��_��~�����u�)��4#I�� '�������(�B��[�� ��		A��w�z~lN��p�J�>W7K'5Ä|B����F2RQ�{�*�>��;!���	l��ǣT�ΰ[�6w��Ep�3` ��g�:N�F�$o����@*�1 t �ק	h�C����32˝M{�=�'E��#咭u�V)�_����:R4�����x8�uӺ�)G���D�ɬ�dt�]=|��y�}d��n,��R(���g�Q<aY>o�e;Kg; 7&��~����̌�.77��~i�v�xt�ӊ����	ab�]^�EmL���S�{�@LBl3���v���P	�͑�������۷>QH�ަR�K§�ЌLM����y�^��#�ߥ\6)�w�:��w��#���V��Q��a��;��a�ξ�s��ʤ�����ֽfvu����g�)����C5�bMN5�͖z܏}.�A������)nUb�+g� 1P���?�i�\�5 �ň����wr�<�Rbw��o-����i�5��)@'���H�E2&�%�����R 	����A�V����Ӡ�/.Q��O#��)unw��H_�(*(*���]�j�]��竃�F��!v�� �����-W���B�EU���x�i}XB�0�5�g�B�̗�,�(	�{�/�7خ��24$I	2eZ�_�b�<}�Vc2.���l)�^wTh���F�1�{}>��"63���q-7,H ��5��/���"7ZYd6�9�R"ʩ�� �]V�د�-c���u���-�'�E�F�嬲������떢ج�q�߿�5���<�����Q�w�-I��w�]�bԃ�q�{����1��y�O�P��!<:r�x}���PXVيPkl�~�l�!��k�ڮ�!-�@�33�lkkk�筸��\�]m2 8�l6f��k�?6�֩k҈�Q��}��5�c��hj7�M׳�a3�j�ΕWlG �R�l1=?3Sl��>T�T��C�C�)��<\d.�V��uֆ;[)+�F䗌"��W����)j`a3��.4����÷9aJ�[!L5�!��\���g�^^�t�_#	�/qju���G��%4Nj/u������I8OI7�:�}���-}�ݵ��PF���沦��1���(?�$&�`����B��J���a��� Cؔ<t�@�C���t�b	>����[
�(�$q�6��cs�H5�[��̰'��()�M@o��f��{���"C����~X�}eL�8���#...==�l�r�rt��؎������X�bȳ��擆mg~�z���9��f��dgǥn�ԥ�:�����;�����g��ش�E����K_����d]�[�j|z�=_79�����7����V�9���M���BV~�5!�9-u�m�uq�Y�6��F�]C������u��o���	��O+��r��kzz�ؔ���<5>�Z�4���h���`����ǖ��s�s����+S�.~ə��tk@z����7:��;�W}I�(�Y�<]�
u\����/�9�p�GUn`xqc,�yְ��7<l�W�-��;���
൴tT�g3rr���0��py�� �ќ6���E�dK�I/*H�)n��#cz
���$�����J�ĳ~	G�J
BBk��d���=F��q��^S���q(.6sb�
��w�Bp7�=F3i��y归��D��(�;KVVb�Po���	D
��:��Z>춲o�bA�T�$����=�l�	��r�#E9@��n��/�H�(�i�3d!�5�y�l/t�9On��z�1��1P����ln绰��9�e��9�=�� Q��w�a�����ѵp�	A�Ўӧ��h����ÿґRQ��&��4D M���]�#��=�	�_?p[�1X���Ae���}�����^7����98��O��Hp����頾j����~ ��0x���㬻�a�M庼y9rN�8��`2y�x���Ծ�lޟ�c!��w33�k�<8,�Q�-mS~aN�e�s8�3n����-=�8p����~	9Vpc���+�Ó��W��E��O��?��H�AV��a��$jv%�T���
�$zy��������hG��u��9�`�&1ɂ��ϸv���*ބ��±'#�R>G1��^^�q'�7k2��}���>7�'�d��@2�P`y����UgGh$Q,LL
1�sP�ʤ�e��267QV1N�m_��3,U4����8 ��\^6����lR]�^]�'�Oq��?k��n�2�`{�:�FY���|�?��0�����'�u�����X�tp�2�1��)���8���x��t�Vq|v�;W��s�`�Z8�ؗ��V��%)h�:&k�n'������̶�%<m1��
s��CR���q������[Z�%��G����5X�/z�?�J��ӁQ��H�)0�;ݕ�E>�u�?��F�|~�}�萖"yV�=�ؓG�<~����R:�Zf{���|b�Zb�zkى����Q�
�Y$��6�r�}s7�fE2�� �����g� B@��{�컦����^-����u�Z��M���n�����p��o�ٰ���k4l�zO��˾EF�� ��ۛ�lb\���ܾ��/}��\cH"|��S�{<���S���Z`J�6�:���t��`�JFJ5F���U�0v-n��Z9ʅbcb[����/�|���s�p��z�ʑ�T����3v�gC�E�m��v��*���#���[���1R�?E�T���2l��1�X��Q]�W��2��{��@���~k�W�-���Q����.�{HrQ
h��j>َ�G���W ~�7,�v?�_G�R�{:�݇EMstű ��j:�k�#3��]��g�|�	{�\�!@C�Jl��o����Yݷ���#E���:�Dx�%HN��MI������TA�R��>�>�[*��ݟF�>������i!EH�O�xMK4"�~dˊ��q����g�������,���aw,�eq��ݦ�+�]�0e��>:� D��H�{_}��n����.RQM�#���:0�m�Ⱦ'a�eTO����Lr>j0?dd��T�� &\���J��z�[u���s��{��oN�S�X���L唗=z���VҰ+������59����j�	Y�� TPI��oT���R r6�i��{�31�lH� Sk��n�1�_�8�a�k���JG�ΔP��1��w>ab>���ћG�=b.@�v�ﻏ��򘓖7K���#>)2�91�߇ i���y]~qd�)Gି��A��Ǔ����=3�AMJUѸ�(1�C��TϾ�΃)j�.x5@��y"��N	_�>_���N���®�Țz��B�� {�iߚ��c �=���	{���  ]�:��s��Qqg�UҼ�c��b��~�/Ggid����5�=��L�ߗ*��]e�*�f*�Ы|�#/�<W)�̾���O�q?y����%ryre��t����ߧQ�&
vdCh��GěS�Ǩ ϩ ��wn�c��Ϸ��l,/??��� ��R�w9��%�="��1]~���;#{蛀�s�A��/�����M���ޑ�^'$ Y���۾/PӮ���v�����v��k�,�ß�-|kY���ǡ�4�,�~DZ�n��!q$t�FI�;�n���)�@�Ѯ�}��>���r�og=��N���� �w�w$�������5P�l5W�U���g���<E-7���7lu��K��X�;"<��=�$%����M�$?��{���(K��#��2
@������e5�4��]q�,P����3�q��$�Z�s��M�;�G�%kzS���GT#1;��;٠�.#����99�ǁy�;:=˭��̻(���Gw��̀P�����m�G�ZC&o������e���d5Ӈ�|��{i���Yau��L*K(L=S��ϸ�!9(���h����L�4�O%ݧ����ɚ���9":X�<��x�w��k�Xv����ކH�ca2H6܃�<�Sc��$do�R&z��\"?��$��u><ت2MG����fo� ����ʃ鐿(�3R�x���'��	�徣B$�`ƪҳJ�ޯ�?������iD�=�D�j��^��0��{6m�1�4��)U�Hӡ �|{�9�@�	�<B.��7}MG��C8�y��m�}�����H�L�Q&�ݑ��I����O����:�����9;��X�d��5����ine��	_�̊ΦL�Y@����ۯE�����[p������T!+vc�9v(GňL'���_(l��]�"B�K�G���i�*)���=~6B˴�#��'V��w��)d�K__�����#iRj��I��f�6�Z	�Q�=�|�c`r��&������L�$�c��A�\+p�T�o���({2��b��zT�^�	��ŧF�1~E�.Ft�t��ά�ꑧ�H����y��}E���}W���o�?��L���F9����i���hup��p9��a��k#��=WQ�ߟ�y�\*��(z�Ȓ��%\)T��Ix�9�lX�Qv��@JU���G�n������u���q�Uu�6)��`�C�P���j�Q�s�ކGw�R������?��x�^<-�G�Q������"c<�\��)ǧ�u� &�u�����	,�0�O�f��}�F�5n����� !a��Y��N4.9���d�WA*���1�j�����#���1�,�{j��/�#��{���⺌G�&rJR*��`B8�
���\&�E��Ȉ����4�.ab_�X��yW?����@�������a+���4B5����(2+�� H�0��mn�oQJ��{��i�����%�~<�ۈ�rjƆ
Mصi��G~;����^��#��E��E��zO�O�|���~6�#V�ĥ
�C�r�_WA����G�r L�)xG���z�q���1	��8��&`\tbGOvh���$2��U�h.�,�럓\'J�o�]��m��e��S�]����h��D}�
o>��H#�K�� �Մd���������/�� ����Dg�Ñ����҉�0Ľ3(����RMYؙ�Oqq�����{�o�I�bQ����6Ot�cs�O����Xi����_��x��'f8Z�&"v�Hmo���$�%Z�a8� Oy"�A��D�'�<� Oy"�A��D�'�<� Oy"�A��D�'��� V;��p"��<�����лQ��1j���~a�.�����N��7�2E '�@����}�ؒCJ\�vo�gF�ē����������v��_ԏA��D�'�<� Oy"�A��D�'�<� Oy"�A��T�|5l�ie)�y5wK<�yf��`�]��}�N�Z��5|>AF��2�Ŀ����X����l��7[�oq�o�5���5e��hs�4�JDT1A�:염pJ_�h�Ry���X�Qb��=yv����NqQ��E�#<�NA�MZ`�3t5�J�w��|j�E�Ҋ2'��c�nk�F�l����[{���8b�����L�0�]񲝢�w�p��\c���P<�|����Z�6���C���9��Q����X�at��^��o��J��wa4:ή�+�=�s_F<MS��0�/M�P�԰ix*�����pTJF��sYV��v�.}㺖��f3����a&�� �{	��{�k�%�����!p����k���1�9���Ll3��> ��D�ag��#��|��H�hm�38�m`ȸ�9���%�uF~������8�d�S���;�{?y��i�<[!��V��`����}�"�Z3�'/�.��۷��ܵ��;���*�����������.ő��� -({�㴺"_�8��С�������!(�9��='3K�L�U(�R���:���[`[Aܚ
���,�9�W!����}-�_g����PQ�=�86�i�!j0�5��2E��u�S�;�@И�B���J�8o���ƥ���l��v���Q��Y^l�����<0n�0������r�f�����CG����Uz��b��u�f'10�|Pv�d�>���Yd��Bȝ	~�?�)�� ��d����T7p�Wd�|tk���x}7 s �x:���� t遬MG5�B?r'�]7�D@	���_��׽���GK>�G]'�����	�����S�d���e��z������\�����p�t(t~�8�	.��_aZ�YnS��������1�N�Un{^M�*�5G������/xi�z"""F"���ngE��e���R�+�>��k�Ou�[�QE��ͯ�\�P�$'�8>)F79U��+Q�ק���PJa���`܆��{��y�S.�����˛艹��{��_2U��aJM���p	B���~/Ȣȱ���E�짵ki�G���I�k&�Q�x:�Db��i���k����H!͛.��̩���(��}�}҄�~��a7 IG��4;���f�[�4��]����D���,���D��<��l�2�t���T���e�=���!�O|���.,��
�����PJaٖ=k��:�`S���~W��P��l��9?ٯ�;�����:�a���u��h*� ����j��;�pўUt���G�cq�����:hR���;T�Rg���c��Fj(k�]���/����.����wX��%�BV��y��>i,�ĦrV4�ʍ�*�fu\	G�O�=�֙����2iu���eAo�L��	��E�?�܏ta�b������q�<�L�����حw���^��z��8�J�+����vԻ���������m.�RS��{�j��+6���������0-uџi�,FZ��=����.�<����h?ki_<y˽�a/`<�罵��䧳�Y���8�t�9&��T�01I���lSt��b�/�J����*)Q�p�[r�Nɣ�q&ؓQ-�z5��� �ƦV��)�]'�>����{%EE�!!!sWV{cU�ƨ��2�&3�\ry������&C�f/Yu�V�sfuk:�U��uo~�uƟ�¿%�W��]gc�=M�t���:v>�aX���ZpFC��T���g��qݎc��0 ��oL�z��+�Ͳ6������#���~ؗ���=M���*�םͭ�����n����ym\\v�Ԝ˿�/Y^��]Nd2|�K8Q9E�d�_�^���|W���lN�̀�|�3
�/Nf	�	�(+PYq�	�㾛����]�cO��?|)C�yC�S,�g�-�\7LPvh=�Z�-U�Isٸ�$�}�mU�k����SU��wb�Lltj��ysw[D`�}�,�Ӆy��o�w'�o��;O75:w�U �4�z�~ݥ�A1f�-s�iOr�悟4�%Q�A�:mZ��c�q����M#w����h��j��O���Sݶ���r�#���yǜ�`���yGtt28�ħ�$��F�F�n�N��D�|�
���w!�D�4�a�!�C��vm���{���}=|��W�����豧P80:}����Ǻ²�]my%�����P���;Lx��x�N�N�ߨ���}a�1�<����g�F_�E��RR�z��T�4V�w�w�"^7�����sGd����c�Ǐ�|�s5�/.>����,�Eŷo�HT�.��JV��wa�R(�]]]�)�w6�^3�n�G32D��n�llmk?�5iť�6��6Hr�����#!����|��e��RF}_nЕ^*HAA��dK��gt�27=~���:�I���� ����zE�%��DFמc�}��"詄�)pmT�@$\��ܡ;*,����ōz�3��n������s����@����S}ձ���O��^?i�A��|��R�ؒ�sTw�
cq�����c����p/��	�����⇎i&&����ʭ��V�Z4wt�W畮��)����U洋�WM���Kfݺ�^\�N�O�����+��iAMͷ�=F�������� ;D��)��Y�ɩ)���9*�����b?O�3���|O�.����i��������~X{�bh���1L�f���^M�`�5ˑ�M|""roR�!���n�*=�����>�I��FJי#�6\��dM=i*��ŵ�b�L��7 l��ȘY����8:u���g�c-�������K�B�=<<��P�~];f�Y�ġ�8'|e�v�ϟ���ڮ�HH4�a\���\4_�,m�X�]�o@��ć�����!�9��%q\���!&��t���n��d�~�P]��Lr�OV�ξ�U�rww����ab��w�U���ySW��2���t�˰Ż�i{�*��A�x�YA[,�|���>}���^N�F��n/�%{y��]3�{t�vO�s����	t�������B�[�u~$�*p� .*$$$E����^C@���ԩ���ȼ��Z"�!W�����P�W���8���pnjj�6��i�o�1 �˶��cc���Ocyq�~¹���[˃��l�L�b�(xf�T���y���2�vR*�-�N������5000�j%5�O���w��htP�oV;�)}J�NX���B���@_a=2�p�	O��q\�D�r�2~ɰw��J��B<��{	�~9+��MM����5�����dM9�3]ܑ���D�n�98:fUzbA�q}��h�k����M��v7"��-33Fddd��ʂ\q%��G�� بY���F����ͭ�AHU����8�(�����9����py%�(s@�3���9[O��RL��z/|O�O�W���!����=��i�*�r�m�Y�4�ǩ�>3o}�~'Q�qz�"�5���Nig��zߦ�NL��v�fg=�?��e@T��6|���
J
*�)�5��tw
"%��ȍH+H�R��1�tw�  ]C� 󜃿������_p�4�9g��ֵ�k��I���?���+�}!J!Q꺙��߳R���u���?BX3�+�+���ɡ�����ň��].~~�W�~��U��<�����`�w�刡$���+F��ޞח~_��G��&�7������q�kтj�&$.i��o�+w�������l�B�/w�=�߼��� Y��b�k.Dc$�����뿑P��J�>9
`0`$��^��,�㵯���b�}	ѧ���@ǀ&��I�O����~��Ni�n��#{�����/��)�{�����{Jп�9�Cfc�222�!u���lGhj��QH��5�v���ؒ�[/��)p��+�]����/�>nWwwsW�1�b-�:H?p���t��AGH�� \��W��I��3GGǄ-�t.<�~?Ҵ7-m�nq�v�^M�&������Ú�xw�Q�S�ѦI��`!�*n�m�7����Ȑ@\x����ŋm�jM�����RH0'�Q��͏�;Ia������U��1A(�H=�arnD�M�r��I��;Q��Ц��4"?~��8����0m1rC�>��HF(�a�DO�	Z��4���1�a�K��xdX�k�W�M�L�~�U��Hm�Ј�i 2����zlz(�'uΛ�f����Ht���.��� �
��ee����#�bB���^�w�D�y��Fھk{S������ґ��8��,JcS?u<J�W�,m��� "�L�׭v�#e�l��c5.�@6�	�r��J�0`��_Y��Y�q���x�
�n�P.��f�kY����C�r��b���h���@�����}&&&�I�٤2{�fٷ��v;�CߴX�n~���H��#��*=�t���Q��x�������;�������R%�)�:�\��oݏh4Q����2F�.E�+_�q|+�Wτmg��6�g�;��=��UȻ�LZ������@iGE<BԻ��EZ�5AM>}�@��Y�X�c%�W���]0��@q�o�C�{50�n�E�Q�
�\��L���Gl��_���B������@�H��>Ƽ.�n.��:�I���Jɘ�+�$-��I،	bƤ�QR�MCr1zW`�[r�����|�xn��Z	�(9Oz]���RCcU����06}6����CՔ����x��`�� �����Ѫ	p๥�����������}iw-A������8�K&:�R�2>>_zM�d�jj���l�p�(��qek+�굛O�"W67��/�@|�LJt<A=Dȿ)��#K�LڣG��s�U>��H?�jg����o�e�y��c�� ����G�O������V���b�
�a�f���ͻ�4A�u�ӎ����~�+>d�ԯP�Ϊ'/w�=�
c��F<y	���X�(��%�����2����/�I4��ܻ�����U��.�a��K�n�J���7�d���f;h��K�c �ѓ�]�4o(	�e�#a��\u ��F4�T��v�{g��}� ��^�BL^���l����7Pӕ��D<��b��K���c>;;��Tj ���H`�kEt�ڔgX�ï?w�ʽN@�1iZ�����&�0y�_[�R����:x�6&f��Nim����`�H��*w���qfzj�$�����4|Ћ=ZwD
��g�@�7�7a+[,�IL�wн�K8FU�Th��O�i7�H�[RRBl�����D�w���&��vԽ�}�/\L��X��Xw���VWW�������tn!>�5\���x�ne�+�tJy��36��#<�u��!���ܡ:y���X~���I�J��k�^�4��O��>e�&j��Rh��l�����7�Nf�1�hkk+V��{�>^����Xmip8�J��(I�m�C�V�po ��@4��J����))�����v��Nf���r���kr� ]��	A`�L���@[������4�0v��% H߹�����Ĝ��x�aWp_� @;�.�Ycե���k�$��G��fff��{���w��}+(�rt��R��T���z����>`��X
�������.�� v���!�io�����؝���{�� ���W�^,��(���j�l�	����Q�g}�h&����Z/Š��9�$�6R��w&Q�/���<A"��ܢ��Ø�X��A�حI+Ow:���h��奌L0�_�t���x���K����@&]EC�C��ۮ��|���W[�W0B�<���;3:�W+�j1��|�xlA'����Ǝ��Y����>6ϭl�ߏxb
b DG��:D��L a���EC�ecxyy!j�D8����5��z��H�k7���{��0��^�63�м[���!9�h`�)~�6u�#G�|�;e:y~Φ,�# ��!浵�\�4L0v`> $NC�W����+Q����O�@o8 �w�6�r�A��z���[Oj��Qc�|n���K�N r��R%�k��#55��:{j���6���T����sMD�Q��ќr�[337�ogH����)i�@���0!�����]��I\�@��/А��i��P;I����n�����(`��J9�����D4^SALWxf}&rϻ�� &��?d���'z���b��RxI�7@Y"�J�#���bK���A��̄����'PO��I�}�~�w{ޛ��? �3�i&�l���ˈIJ
��ANr��:W��I135>{�0���3��}�ѓ��'�1^�L�<H<7`%�ݜ��'!$,�2y��p]�A��wEXع�4�$��B���c��:d����2

�4����L ���G��l�x�� ��7@����Y��m���-���gɬ�6����ё?�ni������b-�0P��c�w��r�e��n�CV�eM]]���������0@(g�W�F�	'IC�2���HyE��5��i��X��s��s�՘3%XU>>Ë�k�|�=�nu(k�:�b���eQF�������.X�i��t���,+��Y���H�ä���RN�_��B2���˨FI))++V���/e�m�{5�3\8⎺�ѼJx�V��:p `��6�{�7�G''���w� <����E�.f�/`��®�7iDk�"��������K�or�+�ø�ڒ�2p b�N%�5���]�5XS(?Q�1��;"�}��1*<�ƕـH�)b����V8cӁ�I�- pg~~���o��`�3�%L��hd�[+u�%�{��RxPw��B�0͋􌳣�b�����X*iJ��7�<��Ub@�c���j�R,1#��P��X$&NB2�}E�zDN�Sͯ�όҝ��ר�3�]�^��-2�7��ek���Q@ �*֠!H���J� r��慅��V�ޙ���#բeN
F�����c��l d ��G���ٱZ�zU�����VD�;g��J�^mm&t��+~�/oc���9ܣ���ʊ��ik4��=��Q$���Bϊ>8�� {*!fv؞�����7"����IINF:.9�p7 ���E[X���e��\f�ǫk�+�X,�`��bc I��O��b
W� b0���I�_�����|K�v�A̓߹� ��a�3֔Jͪ�{�Y.2�8�V��E���������W�?땗��,�7^���Ðf�_�=~�ӛ��E�?�\�RK��(\y��⽂�R͌�WT0~��{�������5[�Gi "�F��&O.�ɫ>&D���>Ĩ��t���0Z�x�.Ӕq�_�鴱+++$�,:��5����˴�%��%�����%ask��	5 [�;,8�����f�4{����Sb��KMMO���I��t��UUUDQ��������ͫ.��
�n��t���ϐ/J�^��Ҵ�`��ѝ��x�		]���U��H���^�U]]�tI�wP?oLM�����A�����yDK���	������]%����lcrP�"򬻂���_dfd�� ,,�}�2��{`pK�T/�0�:�����S��{X5ɗ9)u����m)%��_W��c�@���D��h�>�����5`�O�oGG<yp|��U��� .`�J�9r�`��6ݚg� ,�~Ql�C�G��n-on����n7�����������	kt������W�����X�	��������?^$�����j���!���h	��Ǟ�t-rD�`��Xbr��#WMCI)��=�*�?|k�J�v������N��ń��8׆�āZ�q�=:�����Wq'��]H��C�O� ���9�����?baqV�6�Ǫ?���$`c\\��D�)-7��󫪪���5����ɖ�����U܄��T��:���K�٫ey@�죩i�����+&��X��0L̫�z���\0BM2���r1r���~���C�L�H��oG���Ί:�@�����dK��,�b�9�Gt ��~Ħb��L�D���^�W�)1�u3�m����['�*�c���>����9@�:6�uP���ꮜP����1f�+����}��DY��t�y��;~���� #��ʖ�>�w�K��Hlp�'��E��/>$�+1�뽴<���NϬ�4��I|�e1=���m055U�͌C���x^-w�.���G�6�y�J 1-8�Cw�<����s�73.:%�E��i���Е ���>�bA
�F�U0�&_j"���H���+$�
fԻ�ࢇ?�A���eqX-�;=�>"""Ҏ1�	E�����x!�2�Wl;A�T���3��Y����Y�RRRiJ�2��X�r���_1($| �(�:�Aa*�;c���t��$��wF��`Q���g����&������{IOO_���񱙹�&�*(	!qIz-6�N�x�MW�F�V��� �,@߰Ȥ��9��~��u?����}n>>2� �:��a4aEEE�n���R%�݄�Htʶ�����������l�x��0�=�{zZ �5�?� ��x�J������`
u��pε��(49��L �it�8:;�4�&Df�HC�������� =H:o����?��A�A�A������Ջ��p\�13h���[��6~��Hw���ɛ��*_
t�'���*�\��o1b�E��oD�kt&�?������,��$��f�����~�AՄ���[�Ñ��@�!����x�y�����3j�[����� �x@��v(c�Ç�&v=o_j5%�γ4����_7��x�fwĳ���<�ر��L:t��(*R^�	HI4�O+M�f�]�;���<�[q����}^]]]M���]je��}���8�I\���P�t�
�A� ���]��:�OGp���uc]L�f+�it�>Nӛ����,���;A�h�����3u9�ym�A��.Q�M6���1�����X�O}Á�=�� 
���O,�,�$2�8d��.�-�:cG�r5��X
�n`�*��A��2Z�c^�!isY����d90�Y7�aⲴ9Vb�H���<����m9Zw�	n��چx�$Źg;�XF�3Y#�����zJf��i.Y�,���6ǝ`�C�;��=�;]�r�Y͆�ӆ-��ӆ/��vr���%��
�eyL���x�#�����?�o�����l�~�B\�EA�;\��4m9ç������3�#��xaǃ������Q��(*��0�
_!��l�VG���yf,�z�>�M��OO��|�U�����Ȧ�"��	��ϑ�P�4b;W�����*�@����m�ܧ����h|�m��0�]�hNj7�[�Ǟ_�W�[�up؜,|����!#�!US�y^hXS�����oY�(ذ�F
������5_-���\��_�Ӿ�S%�Py� ��O(���w~�b�h+}tĐ�*� ��c_�� �8z.+N��#�9J�vH��b� ݢU��9��*�<��:�g�Ki�|��c3��S�^	@�tn���x u(��ѻ�
�#����ZA�����lVV�\{;����K�E.n>������.�����'���I�s�Vy�����<�ł*�PQG}�4���b������黡P(�@�[�D�S>�SgW]Z)�o|�jK]V�̘cQ�~HM��_�=��$���(���j�rr�79p:l~���y�O=j�i]�=Gf�+�<�q��G"������^����%jQ�RU*��h�V�@�m��P��}���\�����kȭ��'���qI��h|87�'^vp�͠p����~N!E:���/>�Z-��3�I�޼����̳[۵	�,���^�\Y�9>C=�q�19�y�~4{�f�t?� �r��D%�;��R�^C�
깽7z��P��JGvl5�N:P��b����F�\�)2��O�4f<PY�uxא���Ǯuإif�����|Y��f=?�:�=��:�>�GK�z�$��= ���^�����v���T�ǢvD?[�{��'q'�R��ǱGu��;�v���wO�Y��4_�
D��񋯉�L6���y:�佑`-�Ǉ΂����Pc��Os�//K ������X3�2����br��i�7JT���ʮ����Q�m4��W�zJ��ɰ�d
-{d�X�y�����C<�����-��9�C���Oyr;���9������G�f(`�g0�
�èD�`m��S�{5�_��������A��ق7���xeF�d��C��#ɨܕkw3\Z�OO ���t�-)>�tyl+&��r��j���/�s"�M�b�-Q�n�Sђ��7�`;_�����+aS�(�B3����-�v�=�T�w��y�_���%�V7�n�f�YP��Wr����h&uPx�J��W��f�9jNM�B3p��b|t$h�����Ġ��vsd�ZOO���o��-5�>%F�gaQ�Y_�ݏ����-�z�$�Y��[9h��aP��S�1'D��V�����������`�-�%o�[�?L<K�c�ԷH��G,w���j�^�1(2xxc�������H�۰���N:Χ�N��=\�:N�T�4]g߫o�O�m�*|�����$��'꾍EK����j��{�k�P�4�����c�L��+��$l��7��X�9�[C_��1�rBn����>VІ"��r#5��l��,�����k�őb8�zjo=�N�����7Ț�	�+&��g�-g���0oFg�͙�o�@G�/���)���B�٬k�j)|��?��b;%�AϦ��}B�Wd�3�\�zC�po�)�I���v�*tV�`�ҭ�I�+��JˌM�|p��u	.�v�x�1^�x�q�n'ً��ʓ�9��b�~�K�_Y�e�詝�yB	,�^ܔ�D�H ��5�~�ҠZ�8x:�".}y&Nݘ���v�<x���E@G`��I9�@*�%r�-�62eG��^��� CrãX�&�sG�5Q$��P������/�"���]��t�;������]<p�1!!xee%&6�]&]%���oq�s�m�W�|���(W����6<= ��08�Et�(^j����K���4D��2�z�Z.Ym�C���L49,44�u���[T寮�!����f"E�[Ra�!j[�5����p�P�J�!�S�`߮`@�ڜ+����Ȟ�&�(j�\��G���-}�D�m�x\U���XR������ߙ��Vf$��ը�3X�g�\l
 �����?t��y}�`�܌�a�"��+T2� ?m�m�&BH�=�����A�/�A3Tq����$�,aR���C�988H����M.������hzW��/{p�ٹ|�ܼ�� �X�Q�7��Rh��j6�N�9 65넜I��F������ەEl���Ԣzgh�޴����P3�oj��˲x�+������
	�v��eG&߃E��>�X��L�u�0>���̹b�\��9���N9+N������^ʜ�g�w�9����i$���LGNN�)��t2�u3++V��%H��J��`D����1��	O�~����5Cj1�������1�1��O6�;-���4�ɨ��V��]��}w��w��		]OU�d���6e¡�k<B.u�L���Q�(���@��Plա�+�cG�'��5��̈́�}��3��ML����#�(:nm3z�w�C���Utב��Q�����}�&�}���v8Q�%}���:,�f��'y�����t�33�,/�v�λ���F�ݒP'H���'z��6������&����2b��
h���S�~�Or��w���۝鲪?9��icn���Bso���|�G)/5����.+A󷽴&?�l�F���El����U���|���t݋�o����}�s��W�.U���?~�N���Q�l�A��3�26�n_/y=���m�a������$p�s�8�[���v&7� )֘
T��V-}�.q�so�4�7�<�vf��:�x W�&�D����S|������ݔ�T��PEh`ɖ�)�a߲k���Q��k�W�igTz�QGG�q��g����<�j�ڴ9�����w��1l�=�*��*]�A&s/�R=%��{���n,���|Btj�����H/�a���+�����d!�0���{���8�Kd�c����xu���LE=�\I���?��_mX�9M;b.�0�C;�B�O_>��&�ո����iN'�"1r8R�@{�BV��O1{�N���Դ�qe@���43!���h�ߍ8��'`�4��Ia��P�X��9o����]����d�4{zm��X�r�h]���:=�:w��*9+S�?�D���Za�s��hE�F �ڑ�߾-������,,,<��<n���(;g.d��Tw�]//��u��,0�W̡��jJq�#�|9�\�R֥ n"�&���:�:��H��޴��N@�I����m0����$-��v���*o�##�`�����}\�㝩8� �[3u�w�iĹ�P�|�b���t[��p�o}���A��Ь�B��j�:�d����p��l�AYN��رw��u�Va�O�X
��ɉհ^8�M�4===��� �=1����s�=����e.ך_G8k�)}���sa��A����کZ���j�bՔ�lf0�Wҋ��˾p�F�J�=��YVV60?�(i�ܨ�z\�|�����x tiIËɻ��>9c��+�.����o���v�q���'\�O�F���������ZuAD�Ύ�
�`u~f���%��zb��8W�EV$�*F%5%b1�9s.�C��_�e!���Uh�̕o��t�1�t���mz�~,�P��_j���6������o߾}H��n	$a1>������5��W��h
��)� Q��-�U�wƏV��s�c�޴��7�1LQ�G[%�be_�W
��Y~�T~ʩC���'\�%|��p�2���Mz�xH���IE�0��J�8tbb���E��<��稨��r�����׾k䐔�딼���Γ�����)1�����������3x{/�ίO�(�4[�o<Z�M.�����p���vI	N닅��?w��VW>��S}�˨�>�e�����<�j�~3����o}���;5m$�*��f����jӑFԒa�o�AO�ddd��L��`������> ���hN��NB�y��t�Um�#禮��<�4@a{���7S��͡��䩙!�����T�j�)5b��7�Җ�w͖��l3�����>�n���Zu9mFy9�4!�}�.yf�����xI,K̈(�#������R
u_�ٵ�ص{G?�Q��V�*5���F�O�[P޵�4P1�7����~���@�T�eO� ��Yr��k���$x�G*����V���h�w��ɤ�S�pss�2n��?���ה��D��j�|��m�TLm��V�������/w{�S���U�).�#�{dR��w�*��z���`ϫ�
���ȷ��y��tZ�^��07�ʚP��_%68r�1U2�LqS�D
���+l�ˣ�V�ǋE�#�Rvvvf����8��׶ƀ;ji��Y�(��D�h��֭șMϑ�ӣ��u��;��,��YAM������=D��aV���5$-N��d��X�_ Ap@.Q�r�<��t�_�a~wL�ڠ��ڗ��L��ƈ�zFZ�uU���JJ�G��[�3.ޭ���[�}Y�9�0f��k9I�h�Pl�>L"I��=0��u��򲲁���A��a�G���, �,Wy�wL̚�)�k��#�Pu߹�/�1׿:�[,U1����ᘵ�?�2��������U����L#M.��Y����F`|�S8�g7WM�C Y�e����/�e��:�����&[���ْ��7.�7S�1���w���gGn���x����
���7�G�R܍Wh=�n�aY�[�Ύˮ�ig�gPD���]0`Z���쯹��$'����q�#���,�>����y����fz\_�M���0oKå����_�_���H炵)��;31�$bo}�@p/us�'�ٍ�V���4��m ӧѰ`C��Q����:}�pA�E��
ջi��?�(�t͓����mB#�E��7J�TN�<����z�ӧ/^�X����Z�:Jg�1�0�t��W�0#�{�x�5i988�kT�sH�F'�Q���:�Q���g�.M�Z * ��m��aA�u��Լ\�i��,����
��g+�ʪ�%_~�\:9��æ\��\��)���@�i����[�{�T��v'b���J}2^6���yS�z5��?+hB�DH��F.^>����T�G�P��v�k�k�f��L�3'���y�Ji��6v�ߍtP���������Vpp�������Ƙ���������Ns8;�!�jq�@�K�-k^�u�H-l��h餁��n��@�;��L���W�=�&��H�m����E�,ɰ�c��m��0)���P����=�N�����R��5��� *��@n�ܓK�tJ�YX(�%�`�q(ii��yK7�b�6	��<\�޽3p��׸ɶ<�����)O
�n��\mϙ3�9ў�%&<?�,�}2����.��s9r�z�r��|	A�Mc+&�YU�y|��)����sG?[F�߇Ey3L���n��n�$�?Ǥ��^Ƌi��"��@�G�j��gbc���3˷����M������W5 �����R�Kn���J���"�55���r�[���a�O���q�"�:n+U��쳟�l��X������,���ep�a!:Z��I��Q�3R�U�-���w�Vg�8�ޫi1�`;������;��,C?��`����9��doc�jh���d��n|��{`~~~ ;89؈��~�b�  �҃���@���q����<7����.�~��w���5��?������e=yW.^������d=�\��U��p�~w.P"��׹E2����݊y;D�o���<>����Q��ٸ�w��߃
E��oVO�z�Q�Ɔ���y�p���k-)�*�%p����XXXT�1�%%��_ F���"�)�V�TMz�	�+�<������q���ʕ��{~��J����0j~Qgi}��印	N�OַW(t�@��h$ҿ��@5�U��T>��&l���:ɽ����$]� �⛘4�3Z"��̯����:��q���� ��<V�_N����VW�����o����/ ��}�G��ӭ��D6A���$���:	Ȇ�"��@��~qP'�}�V�:Gr����HCPBg���p%�A2���k'h��V!�ע�=�W��z�^��
d�x�U���N'Y����A��T'�&���n�6pc6;�ef*]N�ɑ���y�,'q6�H8[�WI�vP��O�̱�'Yb�1�
QWW��a1p_InP`������	,ؐ�<0o.k#ygA����bnKCX���WI���M$Eկ��#G��&�K��)�P+\�S�[W.MnL1h؏9�,�G+��Bv%�,؎�l[�-Rc��oTx���֖K!e��x��I��YII��y ����pm��0���e��'1� a[��ɂ��N��P�T�z<�]եf���]�6������G�$�/9�:X��w>�`U�$�f�fJᑹȠ���+�n��"�o��਩�����y$�RX����s���D�3kpa
j�|M�IP;�a�~m97m�OS˩��=>2��q6�0�o4v%�M������x�y��O������]ӧ��rԦ+�:9\����VIp\�F,�z�M@�¢v_��Uh$�)�;�[Z��>����$�+�.[�!�"W�l+w����Ĺ��Vt賑�OSx���U��M'�dCդd�[0���%钣3T��Zs"��5[�7a��^>v����4�S%zp���e�A�DO�OFa�ͩDPR|bRR��"e�ɋ�Q���f~ �>}�$g��zC육;��dPo�|y�GO�9���E�7B��m��^ý<��CP/FC�/y���j� '���C`3��ө�ʹ�,�C���]�&s�Ž�I��`5�*��Z����b��O'���ܜ�M���4mL�RR\\<g��k#dm�)1��\>��}u�Wҷs� s�6�˚����l��'��{�8�nŇ<���P�+ݟ)�����e{���1�+;����P�(��v�8�A��$����V^�	q]*���H�㞈�q�$k�\��9�C{�P¢�=j�:���i���N�V���e���v��ݠ ���%��+:w�)�L-�䔙[���|��3;;��y��G}Ν�F�/V$c��%1�f��e��tG���� �$r�c���'|T�{��5���'J��X�c���DvW��gټɽ	����,)�������9-D�q���! �� �|��j&F3�S�*�c����nߐ������c���W:�:~Ts�I�P��������}9��M��n)+��r�v�{[�0���B�DS���8G�
�C�,X���"���$�z������<)2:~�ݺ
&7s£��0!���t�nnn�jj��|����Ȍ`�ۂ���-� 8�J˘A$&�x� f��r>{���A�-q6���^���97S /���Y/�Kh�vv/Dx'A����=e��Z=c�<YXr�}~�[���h��k僴ݹ�R�(��HlȺ���Z���f/�S�^��^`\S�>�]��`iOFF&���0��FC�,�shԑ?CEl���#[i��g���g�Hg�+y���Z�x9/{n���=�?�m���TYe!A�'9�A�:G�.���kڗ<��=�0>�Y)Z��kCt��T7E����~/���hƂ�h��Γ���+���o�R�y	�/�����М���2�բE�Shvv�V]���+z�����d� ۔>Hj�h�Q��/*��-q������ǿI�ߠ���c����WG`���.\��bn�|5�H��C�Ǐ����W�mz�Ճ?���`M���]�)�R^k�*��6��a��Ͻ�3�^��<v]@�����Q����SN�G"M���B�nӑQ���� ��#�sFdZ;- �Q�y�����6�b�F�\�?B%�C� �Hy`a�ڦj��Myw�s(er��r#	�M.[{�oU7D�#<%�%�C��IfXÌ�ע�^�{�cK���Λլ�bG;Ͻ��$F�%�CF������G�ͫg�F�Cn����w���X�7����O�i�v�%P�6=I���a�tci��Eqo��yLN7��^\+?�y�Ϊ�H�Ѭ�~Y�8BVi��?wZ�c��dS��T�B~>�]�-�OC�gg0�{�t\,>���<�%�Q$��)�=����98��n��[n��o��mc����w�9�kl��Y��w���qzP��8W�:�	|���B 8��l�������)�85�M�2��+ɦ�z�W"���Z��>ϱ̞����47��)�Y�jk�qgt>��cwSc2ԧ|#���= ���ә�X7���}+O���c�S�8>>��TL.��ڨ4��m��<�
��&�,��Na۸;Z4p��������MF��[坭��YFԚhf�%@�J�u��:�΀�\�|�c�c�n丠$YU�e3_Q5*;A��5����ι_�0��b�2��K��{\�n����0$,A�����������DI�(�C1ܪ܊PQH����?IC5���������ڏ��:+[Q.�ν�hfy��Y%d��?S��5���j� 	R��7���M�~��&{��Y�,@��q�!���A���J��2w׃��6%���(nHN�d=P�y�__����V��\��f@VIf�U��2��o.�L���d����
7���ּ-�}J��d�}p�c�E���z�63X��:�Ӧ��~3���������D���pYP�������[AR*S�%����%��D�rKM�:k�?ܛ?��O�7j�[^���;��Z^Pn6b@q.MH1pI�5��ȸ��n��f��a���3�QI��Q��%�e
0р�?}X%+#���B�c����IЄ�B�+��Y$P��� ��4F�m,��>R2.�����O2h��4����i�LQ)^�f=�wL6�����fD)GJdw����9z|�6Eml�2Iy�����dqs�����3'������E�A���p���>�z�D.�\�T\L�?_�P�x���H��ڝn���o|dh$��7����QN� �{Ѷ�i��z�B��21�[V]�ثfI��n�ދ9��=�-Ā�)���x� Bt��"�?��Rz����ƓS�2x߇�T�K�������a�ׯ_L`��-���+�B,���~0�ٯ���a@�v�{�'�\g$���ڟx���#f1Y�;��N��0CFL�XX� ���� +U����ء��9`1�yh\u���\�fG>�\�%�3��c�=.�̬������-1�ߥ�G���ߎXH��G���b�r�t���E'�5 �7�ؤ���DF�sY�V��ܗ�w���L��ȃ�j�>Alll��ǹ;:;uK��r4�e�U�wF#��o�����������-i�m2�nM��4��!���:��yO�}��VmD@:OMX�bf�m�_i����������)��n=�Zd5���Z��ͥ�ٯ�����C*JY[[���A.�LY�:%o�*v3���g'��X�Cu�졀�d�^�2��9�m������ �܌��zO�M���A�ק^���϶g��R9��3�I�CBB�Wnfɦ��U�{�
8�6%NDmO{�E^^�Ł�T���y�N��Q7Xb�H�d���@�π�thD���^�N?@7�M��)g���J��<��Q[kB@�[Ȟ\���H�q�L�;�>V9�F�&�B��	�f�b[���t|p�ȅ&�ѥ�\��b�}���:qXj9=��=��K�]�ف������k`�}��`�"�hx@]�b�Wh7�h}�&Mdp�	I#W���{Iޤ�Yg�A�j��F�$L��q�n�d���\6:	[	�D�8��i7}��+�9\���?#��A����ϝv�Q}��V���:��� U �u��0
O!'�->B4�5߭���ț��n{e�j�:H�-Ԏ��7Z�j�$j5�3�Q� �S<��XF3���c&��b��$��B��I�b�x�5��1� �V@4%W��O7��D��/�� ��nlD2*���)))�
B�G���9��T.V�vvwa������V#(Wf&�~�b祓��CC�HkN⺴�b���h�5�� n�"�!��ݑ����45!�Ak7a� �hɅu�`�-�*k�/������C�M�D�OwFs����>b|��2�E���dx������u�+�Rq/u�MS�_�����1���Z+��-���n.�<��0�X�@�����1�}���C��TJ�����b�Q�+k��1�=�FH��vn�5n��D�'������PRS�@|׷`DYYٜI��׷ЉP�e���������[�!5aa΢L'{�܍M�_H��.n�1���^���T @��7��uٓ�ho@�|:�.S�G��f4���[�|uCMe����������V�l�վ���>B���hSsyՙ��ׯ= K8AQl��,I�����&��m�ɼ���~��n��l�^��B~�[vF6n���Y��a2���2��gגo�4��N���T�쑻�:�ݚ{hҊ�B���\I���8�C�u��Ό+���-�Q��M�Ca>0�W�/#�t	�yF��z+�����r���w�?��Y��SÖ���.5��}Y�@ؑ��I��{i�ƪ^r
C��yxxh�X�]��	�\%���"�l�k��E ��Ξ���!Gr�:�
����0�|磹�HK��U����$���>l���ޝ2�o��w'���b^2T�b������ߋ���\�1^���9�$���ȏ:\j�\'}��Y��4j �2����ď�b�� ,����l�e$�U��0^&��˃�l���g5����l;�j=�����0��x��vܧ3��(�h�������Wx��Ux�`V`~������f�%?H�\4�;��f�2��w�hZr�l���_��7p���)��S��<?�濥�G��Q�(��:oC�a5�Nz>>�T$�4N^�[�ͪK�$��2�\�q��$�]~����2ԫ�����ͻfC՛���z�e����dm�>�>�~h�!�FaLtc�L�s�{_\}?,��j�[��]�Ƶ�M�=	�6���b�L؍]>$I,K�
7���TPPHui����n_i��O����� �P}��7��c�m6�z搂+�=11*�)��B6����zpd�=�`n�a����#�f/��ET��py��7iڽ�#Lq:H�=^��T{յK#JSVV֭3Hw�|.?[#��WwEJv��������믣4�M�[��]���z@̛���K:c$����#Jh�Lh({���x�����1�6��/̖�i��H��
�@.l�&�>�ɳo(<ǧ�<k6���:�B��w]�,��,̞ɵZɵ���fQ�U��]�f�gǓ �Ϣ�`	Ȳ�����:Ma�	��)���>LhB@���I�Ď3(�W��x����'��KO6�+��Fw��z�,���QJ	�g��q���Ϛi��N�N�&�kG��s�>\���y'e]]]�G5ݰSj;x%Ҹ�׍��C�$����D�K� Ɩױ���BdQs�n��������({Y�4Brn�r�S�H�7@�������2�5�������4�v�aA$9�C�s>q;�&�s	"=o�o�����'Ot.��S~����5k�T�R0�zHL����T�K.n�@������ ,x����r]�b
%L=wP�\�������Rv�P1����	v��\,�aȲD�����~i�|i�5M;���l��{�3� ��c�
���`ێX홿;2n��ܶ)6����>��\ZXh�!5MH���k��o7��C�g_�EZAZOBDK�0�X!��ɪo�jܪY��%�F[[��*�'������hhhdhrt�\��%,��������n�ø�
���m��������|� ��/W��w�,�I����1<=������0���S�**�Wt��|b��W�/�&k)�&�OĎ{��燒���*"��c��|��*�7%A��D������_��~f��
�u���e�^������q�_S�u��и�}6�<�Q�7 ���<�L���w���5V���{��Sƃ��֛��X{�&�>~�>�PZABD�.EJF	H�� �9�Y()�!�膑<8���1@Fw7�.<��O�C��u�5�}��O�{�]}F�3@�8L���ѭ.�R�;�����ſ��>�
z4$r���(#��Ed����D?_Ƚ�9�jנ���k]��
``�=��4�>� ah:�(�ӻ{#84�kZ����5`��Qm�y}V��R5���^sV��&B���\�~z"��G�@�
��5%B!�Q���LMO"Qn����B�y�����K��TR��>�C�E`ǉض��-2XY����D��b�����Z��8�$�[z��_�g�E��^��[X`_s�# ���4�f��X&n~��~}M��GBǎM��ԭ���_X�R)����HN)�iWN�E�L���`�"����5�2�jiP�(ŕ���c��� ��DG˝��Ua78"ڇY������e!���ƽR7t��
���� Fqg�T���k�L���+d 5��D�d�x�z�Dy}�S�:��6P�]Es#�Uyj��x�R��1\0��mX�ѝwN����5ʖ�f6�4����������2
�6�rX;az���������	/�:�R��iػWF���t|����e���"���dffU� ��}N�]�jf�*1��RG]ȳ�{�'��oڰ�)Q: �n$x�+��Yٴ��ne	L:$��/V�샟�����g֏������=M�����d}5޸�jY08������9�'P���-9l7�.K��w���0%y� ~���u�2��F����*z�H}(��d����C��886����G�X����JYg��D657wљ�2��#!*,��DK?/�Ժ�ùƋg�`	�3"��؍�Q��Uf���V�+��ʚr�1��ݡp0��ӗ�c�L�FT�9ҟ��%�,����y9���C/�u6��žEŷ_�xv�?���y߾�A9�i��Ωq,����n�v�Gk���D����	�����׻��]�6����R�cVTU����O4r+�9V����P!�ߏ[7���Fó�n�}�S�-��"�R-��:):�((*�Q=�" �aV�U��ܲT��A;XZu�ʹ��w��$8�^Ç�_5TU�?�<�0�^5���l4U��G����/.֏=<�]s8��D'�8Ȃ�W�^J4����4�{ϗ��O��w#�jN3S�q��]�U�P���A��\�OP�����%�CE�]�+�fK㻽�Q@�#*�L�GO?&(כ�{�dSH��	l8=8���ܕ"#c�"ݐ�t�`�Р��YB�g�����%��1��'�~�Dm�x+���>����@e��6��j���*���Ǚ晽]�y� �
�.'��M �ڴ*{舘{��~�����lhR�މ�S�KJjʆ>i����`F ���/l����$�����F��l����	n��i�m�+RBBT���~ݥ�.��+#�!%i��q"W�/�hw��S(��.��;l����7����!�LP��]�"K�:XȾ������`�R��#�t\	��;Q�6���T�r�>e{�҄����6;���:�ГNA�-��״�;�z$ŷ�BVy��eD�4�Ud�7����X��Q���V��:g�l+J�4���V�������/� ֎�Q���������<ƅ��/���Z���*��@fy0��������&E	�����Ŀ�뎶QD2�x�sD�3��]����4�O�t��X3�d���yN�EG^d�є��.��_Xx�Ӳ��6�ܲB�u�[�[h#$.������O�y숢���P�ylA�C�ŉ���Y��`���GB���4 z�[�l��5�J5�5�����e��+*�,�r��'��ݟ�*�ߍ��/�O�'o�������<A����_H}\ڿ�|��~gR���/�����#UU�`h�1�@S�p>v������j�=�E��ϳ��Tv��m}xL�ĹΤD�.���_��u`j�$���
�܅��1Q0A����*XH���J��l	�r��"՞h���]���w#(o���t4�1_��Ǵq�Y�L�ooN�(
3�� ��|����F�%���Ja�R^��_�*���*�Y��a�|�9y��4�+����`�ʏ��ꥭ�Jqk��o�/V�)i�����`r����y�qE�>M70k*b��;������k���4_��s|d&\�_3��Z0�Q=_�c�);$��)����$#Ż,���;����
���1O%E$��ՏP�8��{\�;��t>�0S�3]RL�Ϝ����R�C�U�������#c,�j���*�>>�ԅ�|���*�7�cf�ӻ0�6�������}�@b��x�����B���'�3���j�W;T[�*�ei�f�[�-�\:�	Q`~ˏXsy�����!�D?��bL9fjK���=�('�\�7|Ǌ�&\NoSk�	�y�k�r�n�Jr���\l_�F�È�2:XW��G��dL��`�q{�J;��:S8�>\`��Zы6�%��;�݌.N�NxcU����J~���C[���-K�;*v*v��ļ{��MZ��!�Ġ��X^V��Z��<뽬o���ݫ��\'=��ȯ���ϗe�,Wu��*!v�12��w�>���kI���z^��M`ۿ?�(ﷴ^E�Y�D���|ޅ����ҵ/D�:�U�}wiX%jv!q?Ȏ���c�������R�!���\n[�[�ֻ)�c_�Z,h,��Ϭ���G�|��v�\�V��^-6����IE�Zl~ܝ���r[��i���=N�Hr���u�^��
�;����|hy�\�/������oa�m��C�+}i8'.	��R�A�Jje�(R�mE:��w� �R�o���콺)�����$���:T5�\�xq;���\�/˽�������#��-��f�RWFE��z̽q�Z[�����e@������3�&��O���ߧ�Ȯ,"X�\��m�<�:�-� 5��<��X��������M�.7x,Di���{.9yM�_�A4����0�=��
���w�Wun���)�
6v?%�Žu��}��<����+�2��R�=&�6�&�yǾ���_�Ҥ�3��ZA�U[��]Ǹ� SI�/bo�{�f����}��n�)�eޫ_&��d�Z-��{^;Z#MW��^v`\:E��q��Ҭ�]�O_�z�Fʗ����C3W ��?1�w���b��`�lmm�,[� M1�ʘ����d��;^�)ι���W{\��В�ZֹN�w5 ˹Wu#W� �N���D�)S� ꭏ�SZ�zM�ձ~���I����&����6s0��w�e�����*�bC�m5��b��ư���[OU�u�1H���|5�Y��&�<��w���ݴ<�8r�z���ȬRiR	��ڵ�m}e�c��7h �B6nΠ^��kdTϋ�8�.��}�nâ��ūdWCxQ��O-���e�֜M�8��@���
����D(w<=x�ܖnO�9P�M.����_'X��-����� ����6ɑ[t+��W��ڼϲ��ձ���:n	��yONa�_+��s��<�oXr����$�{q�5~��S�^��|)J��z�a���v�[b%���/��w�X#D�ww��e�Hz��3���i�3�T�*f{�p�{ؒ;�J�ɖ���S�	�e�E���ݚ��6�H�V�W���y���*��<Bz?;`��uQ
jO�(�̶HNOg+�	����vU���xzj ��f'�l�z�U`T��?\$
n-RG?p�w7�@P���ӽq'5�!l��%�}�����.�eoh�H=��Q�d*�)5�K�s�օ~))����8l�4�E��DjۯY���F9Cj��������Y�eBN�;�mAJC����4���lL���k�]0F��T8B��{ug���{��Z�xz��	lt�U��^��_L�0\­i��e!�#�	5L��ɕ��ɩ=�򾐱���.��k^��Ag9 1��\e2Q~PZY�}�5b��22�s�i�u�>gN@Ί}W���i����c4d륓����ܖ�Z�Ӧ4?���ͻ��h���� WP���\�g�'��bF���׊
9��%�}��_rKoO��H���C��S0�Wr�E�m�`zC����ȍ9H-��L�x��t��u6<�1���\�W7|D�Z�ؔj_:<�9��@g�q �O&ظC�v��N�g]��IQ3�]�}1������ �8��h������e�(Q�f �"g������*i̘��o��R�Klv��z���Ĺ�i6ƹ3s�Ub��#Ϸf����\�q�ON8��
7�L��u'vq��5����Xr�F�7]~C<����!MeE�Xu���W����s���X�k���P���̺D{+��]�l�s��3�{�5�%&d�/n�)�C�G�4S��6	W�XYl0��ؽoSVZ���ӉY�В�w3' !!� ڃ��"�m�Ҁ�iv�*!����nwJĢ�\l\��o�:�oM�C���B|�������>�;��Vh���[d:��#_� �2��¢�����>D���*��B666?uu>ʔ_4���+Ί~����Ƌ�L������>����.(r|��χ�<����nT�KI�f�B��kN>8���%�}�oX�X�-h�s��PH�c&H��9�ɦ�ֺ^����d��`���9Iv�������U�td~��<�s����xN��gV�N�g�tR��\�F�I�XCi�ֳ��\��Ҧ�|�%~���<���#�u^���dI�]��NXC��|Z;��4�j����-���������?;�w������y��$�n���<-ۆ���m�K����o�2�������&�mXh��K����`6 c�u�!a��S6'~�P�?$���O�; ���P�~i�u�	��� �	 {���uJ����
�ů|dadcQ����>��>��;�K�oh\Yt�RbωB�j�O7�p])�|�u���q��~�v^�MъF� ��R����N4d.A�i��\�r�ٍ.���ƅCM�M��ǣ�X���v���~o����76#�NVVV��D��7�`cd3�^mыo߆�ЇIii��n����_�Srr�"�EFN���'� �B�233�n�L��	No�����\{~�h<��ǯ�t�Kߟ�r��S�eD�h����r	S�0�wk�?Rn|����Af��p�Puvv����\���			I�����������k5X�Gf�����bT�}�E�������$��%}�� =G��(�U��RZ�x���P�x�9�r�=K �m%�� �P��F48ajjj{S�___�����C�q��V���!<���-п`�1�������O��O�	����k��}�$�����̬,�r�E??��z�#3~P0;ê�'J�d	�}7yn�S#��y}/����ఞx��@���e�e�j�����0��R�uQN������=��h�x���jC�h^f-!���#�'�����f*d�a�==�-{�@CW�(�kw�I��	�Dvtw�	�ek���G�.��`)�MO�6����5@��n1�Cc%l�H���g3[BFF�.��C�JS����������Oxv���Cg�\��~�N�S��5q}���T��o�{{������X�yM!�|�6�`S��� !�2�ܘ2��������%Y1ɝ���;al�sU�W:1Z�M ���Ȃ�s��2���}G˥+���N�X�9�=�L(��.,.���r��=z}55r�ʅ_�0F3K����UU���G�z���ҿ��sC���(���i�MO�g��g�-�(Aϋ����kb�����K5�n����I��s5I��㎉�u���F���BX��XH�2rsoG����1�� ��)9�I��5Pꦺ�����ϖ�\r5�K{�Cn�}_�q��m�2:}�{�i�a3Op����kV��4ӖD����&L�sssk����K�<��˺p���T��v?�i9J�:����z���])U{�Uʘ����k�^S�ȵL����oh�����J����H�a����'� e��q�a0t:��x��h3�����i#�1z�"=��*
��p0�Ȏc��u���u���պ��?.u�,aE�r��Viq�x�iyR��-?��W�D}zj����+�&[��R�f	�v�λ�Ɋh'��<^��+%�bƳ���u��������<�l���R��3��}Y��O����Vƪ"��.OF���)�Z�����-w�<��`�?>��-��a��赝f�Z���':d��w��5�Fэ6�f��PNg��Ǐ_
/�=88h�6�����Eƻ�3��.����Ф��	��#�C����{y��US����4SH���k�WV�a����9*��G���e�m֓)�Z���+�Co	�6Ο���Hz(�q ż�]j�<�_��0���Њ�w����T��T�v�����|x���5��vw���wc�F���	,�B����l�RSSUTT�I�e^ ���@r�`:V�V<�~O�8Y�
�v8�pdA��o��Mg����D��n��sm|z�CJU��ZZ���(�nM�4Z�Ga�a��S���KY�����$j@e}�޽��{��.U&w�� U�u�d
�Α�����?8���զ��6�'
�s���:�?�J�~7h۪���8���yy���ٲ�O)Y�%6
p.��s;��y7I�ܮ�><(��ގ�~�%��RǱ�X뫴֒�M�@����{}�|G3'w�lߓ�S��c�`�	�c[�w7����<p�s��G�%�����h���,�, m_0��� (t��wo��K;��a�~�ﴈ\3��� STQl]� _s���&�u�6�0�r������f��`�`gL�wu�9�%,v8�-��K&�k��x/}��܃�7���%������4�O`JOP�O��/''�������(fP��r555�!B@P�2z�aJ����v~��z9Y� ��F|�w'f�����Y�)v�[l뜤�3}�Q��k�8�cq;>8:b���%~���	���- �I�`u���Ut�\2��f�`l�77�Z�:��� 2�	?�;n'���'gd���j��dDCLdl�{%ld��q�l� ��C0vvE6i���:5�ƾ����t�w�m.v���2��֝:_����fh$P�+ic_[0�s6P9Ԝ~d��U����)��3�E�QF�3���B��y���w:S�K�����(Q�M۴oY���k��F�|�(��@SR��?\;j���T�խ�d�q�(Zھ��oj!S�!I�܃g!}����ԥ�7�hR���d�P���H�L�"YR��|8������F=��H2�[;����O�l�o7�|����e��7�2�
x��}F	��ƺO))`�GV�26~P*i�?r��R��b_��w�nf�ź�+*�	IT*V+);�VH~����J�"�%�����6<�(�^B��� =��+�e�J>�n t�E��1f::�^VN��m��.T�S˟RT��u
�d��~��%�2;��˙�EU���C c�^�B��OKk�Έ�-�nD���φ��c�!�� _��~Ei,�[����۬)�D �^m�ڛ�Ӱ!�imO����PUUuQ��DaxrW����g��!}��2������ӾѴK)`�Qɰq��[��e�l�_�C�[���#�뵾�|��0�+C��t����e������O�ҒӚ���|��n��U�o�Fmق)<z������_����#8���6�U��sW�,J�׾R7�[c*��EFDHKII��|S��h*w0n�TQW�@�Pn����^3�������[X;LMt+���J��G`�8t-ޙ��H��6���X�r��zlqd)�͏���R;�_�3��qX0"kE��j��������g�D;��AF�k�tE��>2���[@[�WO��J��������;���#��<%%%� ���ŕY�89���4���7
!$D��d�$�?Et��+�Sʵ�n#LK�@�b�E/�u�����IJ�j|�I�ʍn�hH�6E5s������8W��X#������ONd�V�aZ�lO�-*)g�U��qa�%��E�������&�f���~%�'�A�J�Ya�d�w�[�+���n߂%$$���l�7���N���̬�q���y�\�e�58'6IX�ch2��-�g�:'�Y�<����x���s�ba����,`�Tյ�.�5s|�!Xb%�7�@�Ψ�+䐥mS5�Zx����Jj(Vd�SY^	}6�h8�I�-�����P{�5�y�?���}�Ǌx���qUG�LI�6�귳6%��y�	�Q$�J�j�Avdx����������@M������^���M���V4�J���F�bn�J��-YN�-��Sw
A�ʳ3�2�����g��cP
�F�R�j;;��i22�=}�ѷt�����Nn�����/��x���(.$FG| �����{`�t��u�,�ѭ�%����q�ߊ ��(��M�� �R�EK���u�=@�)G���_3'<}VEB���Gp��Ë�ss�z�مZ�(��l�[�KRb�Ѓ=1UM�M�2�/"���v>�X�tmnj�1ٓa%əP��PPfb��)�_���F�	�輦V�7��>H�6�\�W��#n}x���m���3�#���4���*�3I���C8�#���!���v��)�=@!��"�"�[�!y�9d%�����w�����pO��e�f�P9�������.R���Ǹ7��N����װV�-5w�ƪ�V��@�U\K�Kt�J�9Y�yGz�2Z������;׍��j���2������Cev���`/���;T̪::4===����΂� ��q03��6^�~�z�'F��o�ߪ�w
 :eۄpJKEI9;�����ܓ\g��͐�����%bqcf��Ol5WE��6޾Z������AŞ�J�CuX_Iq��@-G���z?3����|��?�����n`�>�>4���m��y���o�GL�[y�� ȫ�.�� ��Ʒf@�=�� ��N_�]�[%nrb�l�Xw}�s^U�b�x/ſ"�󵸛��� ��Ȧ�g�)n`�l�J~�b�׵|b���Y��q_U��r*��sn�b6�CӒA&��t0��`8PY�=�2��L��t�U?��b�wБ�18#ܗ�[	�hՅ�C����L�W&��,� 17�[�I�Η�����*G� �t/:�E�A��׬�qʶ�l�D�6��Z�3;J���U�ϓq�����tRa՝Y����)@�+���%�]M	����@��W��a0Qrm��:���8`�d���285 �o�V8́V�����)_,��\��PuF�L����F�Ws�i���Rnex��x�\�P�7��@�2�B�� ���>d�w�TX��~ĂK":�5n(���^�i9{=���!2�F\s�u���u=�Jѕ�����=ΑfQ��_&mJ�����Ф=*�"6��vޛ~s����GR��(z1e-�W��G�e��f�B��G�G�3]i���Sm~����B�bll\\Z:�6.DffmX]]�S�"avdT}�t��������V�g�tG.	�sZEZ�VXn��6*���D<���8?0��7M��,a���ћ�f��v��{��끨�;�V�4���mjS���l���4S�
��j�-��]���4���p�D�Bf�*�a
�6�h��=1�16� ��:��)4��tDh���n�T����G|y;�葼���-���ᄚ���ƀ1Ͳ,$Qr��!lFĂI��k˨���mll�Y(��QPP���]�}���;��0C��
�0��#r&�7����F�'7�j���z�R��x���0�
��c�*�6�Y�{��2���/vI�D��-��p��KZ$���QE��!�Z��I�is��;�����K���5�9�< ��8Mؙ��|r�0���)
咀��H�f��o�U����G�����"�ȁ��Q�� �xN����#` 1�Pw﵂Ø�X�������C��ylT�Ճ�ZI��}�C�}-�o�c~�8���/��9��O��4�<�ߧ�6<!K�ħ��d6�p�-��z�+�m�ۮ��O��8���U׏2�`\�]�jOL|LظN���Okkk���&�����H�'���� ]�ܤ<,g� V*����Ӌ'�(�:��ܱ�T�c��ۇ[`��v��P������}䷆��mz�ЃI�+�;��2^�������xψm�*�3#6,9��%tҔ�����Q����������E�j��DC�h�mQ1��5q�����������R*a0"�Ԝl��@�ƹ!&��������z� A�A�Ȥ�x�&��{�#�C���65�G�e][�wdU+��J{�
�0�8+���Pc�w�AO΋e�^���~�[�������C����K/��*
%��n�l���Ym|��yM��[n�������b{�{̨���횥���N�3�rԇG�t���&�� ��o��?iY�-��)*�t�)Ƌ��9߭��;�c�{�A�z�#��a�����'�q�sg?>^'V�L�	����рiȪ9���
��-!��`��0���h�)�"�EH^��X�@�QQQ!��ySs��.D�u��6zg`xްrV�e��')��+�b�i��@q�5�� ����ݻk�n�7ֆV%m���|U����9�<|"�ೳ\��(�JCá]wk�<݈����);����H`�\������4x� �Ot~���Π�ړ�z;2��Fo��U��ڪ�i�<�w#c�+�%e[l��k�����]��ŝ
-�*����H�H������y���U�$ٗ�\��\`�%��?�,8#7���3�N�����𕷍���eA�� ��F�Yn�\�t�b�[C��~ޣKgB�ɺ�FGq�e���*��J�w���j�N�>g�������i)�����\R/и���k����r36|7ц��λ�����5�"�t��+c0 �eeeU�2z�:/Ϧ��������Ѵ��&���_x��{{z����/�}&5��E!��@����r��&���g�}q�ʵ=���S��S����H��n>�u���"�#��7�0� �u��WF����U�.\C����62�5�^��9z9*�+8����rF_f�Ɛn�Â�p$RT[G����t ��������c���������s������IoN������#ԤLG�� �263��'��@by�/���4��=�����{��Նn�Ud���+**����?^�z�z�:��nC�[7����(�I�ɷp�qY�<H���t����=��(mT�01�c���b.��ѽ��/����8T�\������D@�;�G������ 2MO�F��/�����75uu);;;��EYe�> ;{;g�J���n�"�P�R&�&j	�V��U����-�k�q����Jݑ�u�ʡJ<��oG�c�_���@�I�K��͡��<��mB�ٯ�O�u�Z�Y��_�#�Ä�A'�O�bh~�ٝhٶ���4�2���:;/�^b	�k�455� H�w���)۬5�^�ٛ�����R��H#�0Pd���кA)
��j�8�=��g%_�}��Z|B�p?Qu�-����]/�[نk�2�6DV#�a�a�7�H��A��m�|Ck�c%��~gDX<o!���n]���5t�@�.����� �@'^�����ZE�Sb{�gBQ`���A���;VV)4��BՒ��.����C���V��g
|ߥ(�i��#�"Z]z��ģF����U���7pW}�'������6v�Nސ���k��;ϱ��#֦wt��#?;{��H��h'����93��G|��7J���:�)��%��G�Lc����̦,0߀�;.g;AFl�`n����tq���)@B��z?a�Y餪*���*�Lee���;�� F.�	�������)��xa�dF�� �����W��ϓ�dv�ӳ�:��J<4;���Ѡ{����~�Y�T��k�TvGx��̃)�m#�FZW<�v�6��M��UiX7_���
��o�̶�I<��S[�P����#�{3�/�j�?1��y��	w�;
����]i�j����`��>wT��<���!-Y��ViUծ�"��C��H������c���Qb����Ȼ798�>I,N���T�bb���=��¦�Qt6�{
^<ƃ����i|_#rt�6&{
r�0�Zv�����8�����Np7�K����f�W�x9��1x�ٵ��=t@��H$F�����얯f,���p�Ȅ�������A���_�j�B��������������T|u'dnz/�1�t��;W�@�ā(��>��5h�TRQ�S-��Cퟃ��F�g
�n�)K`ho,.uj���K}�J��klb%mi��3�����OU��vr�{54����0J���N��{��{�l2؀ŀ�z���cV��T���RῬ *X4���=�f>���	~c���'  �cx8A8t�sě�9Rՙ�vvn��Ka��!�4nI/!�7X�l�Ay��?QU�{��`i��ܾ((r��/	����F}8X�m��7��Hv���R�n�Vn9�_�=,!fff`V`���qN$ ��3��Cu��k�Z����Ͷ]t�k���7n\�۹l��ʈeH���K#5rM�������J���1��~'��y�tOUo������ݫ���}B(a�)��*_l �\30<L�5�E��"��Cgr$�k����,��@I2Q�t��w/���&]}p���L0�1kׯ�j�]Q��0�1��R��ri@,s�I�F�[�(!S��Bl��L^����~jgMU�����/���<��e��d]Ngk�<RnY|y��%Dͳ�:a�ѻ�4�ݙ�=L�R����b���F�|�t�;�	���+�*��%f9Y�t�1t��bKH����rK����R\R"���R.exA��<��;��p�ҕ��ݍ9��+��((ˆ9A ��Ii��G��]�1�)�&����!�Q��!�ݞ4Q�O0��ZQܶy�,՛�ȅ+1�tq���h��y�=D"z�i��$��@�K��uW�r�F��"BZ�2�';QgH��	���b#��e�ۣ��f7�~G�f�~]�Z���FJI��w����CVмv���������.0\�A�B.�1�����B.Donn���w@ؔ3~|`�Cb��PWn�����G�W'[?%�\L/J�z_Vwŏc�lx��0_u6��oek_����/�1��χ��D�H]��5DB�
��t�Y	N��0 �o� &�oD3a��(�}��M�|�''gyQy�`o���«��IE���z+�^TD(�)��������CՂ`�i'P|7�9�n/�_��m��r�]�]d7JEF�$i�3_t�v����p��{Go/��� ��W~4�u9I�g� �x�̨M��9Ҫ�}���g1B�w�"/`Ȁ�Ҷ�ЈĻ|�Kp-\�*�	�,_�V�ǳk��3��.ҦЩ��J�?K=��I��w����M?Q<+�}��������U��9�a����,��}E0Ϻ�#�j����u�zZ���Y`��Ք��;��-��j������eޙ�=	E=\~�����Ȼ@vp����B�_Z[[�_=���BTA��j�� ��a�N*Z���[�=� ,�c�2Q=�*���!���h���(&&&hT`UChw�atuu����+�_/r�%�,3Um��~��\6�ې����A8K=q��������x��G3��u�P ��.��= φY�dos�K�ǀ>�$�
�7�uS.��c�)QH�e�R�sɌ�����/)q �?�~WзS��b��ۘ�����x�4@�5?�&�������L�ͥ���� !�
�P�wi<q�^�7�hKo�AM3�͛7� �Ǹ�?��J���B
�������G�%�.�-��	�	�C����z|���:E��������Kd�/ӳ�� �PNNn�W������|��z 6����O��,&6��q��]���3�������
�39d�v�I�o1N�ۋ�}��*����`�FH�Ŷ}�Z�/������J_gd3avǷH��x����|��k���G5�F �b��htJJ
X"[/��-�a�'�w���Y󖥞���̛Y��:/���8��m��u�6 ��e锘����ϗ��7d�����}EH����O+�BAY��:#k��<�_�ēu�XnC��5�w���5\4-��/����z[2�T�77�J¤ȷ(e�l?F�����ȱ�G`Ls�  H�^�c�*#���i]���+�-/������}�>�[4�����ǻ���P�c�.͉����ted�W��D�ڈ���ӮzG�U ��8\��x�������CrW,`c^/wN(%��Np!��^���5�k�������@�[����Wߕ�O���V�@t�JY�7=T�pD������=��Q�	O�Ro	��c�2h.$g&o�ۊ�c�g�w0%�?��'���oD�b��e{�.2�n=�Xy�r4����P��_��H8L�='���׉t������,�d[<��$�}�����{�(h�|5����p����~Q<V�ݭ�~�k��n�c���2ZrZM��;���5ܟ���;7��v�����c4��/��Փ��W�a`���[�mv�X/��b;�e�A�Ò[4YHUt�M�����2�Q�{��_��*
�{�F��%V�ڞ�<��gg�G�B�V���"�k,�Ebܵ���al�\�qo_-�]��*�T��ޠ�'c��--�A{B��-�m�Aqb��{Lc�	��W%G�[�+�gY:S�a6z�>�vLF�X�3V�H�OsO;��#�f!N�T2�Nd���IΪ��CX�p�{v�q;�{d,�k�-Y��>(Vl~vU�/9IRZ�����m��l���w<c�(��#rZ6 ��^��D
+�O����(��
��<v��\P}��M�CHЈ�΂,�_kf�����
�������&6�f�"F6%��&Q��#XM	тiu���d����:���OD�ˑ�$a��������1���E�n_ ;�y`m���DW�i�͛ڔ�U��X�c��<C��>x$�3k�;g�����8���P�
�^�1˵I�Mn���pλ�������"Mޫ�zi{�� `�z�[��j��0�`ʝ�H	!�t��E�"ۿF��<V3�t��� g�����;d]ܜ�2�?��2n��2[sӪ�v�����lfn&�՘O�����IԲ�>��R�[ak��.��su�W(4p*�m��CH���G�*�).�/u��BE,�"!K1>o��gfV���\�Φopn�`��ux$���/����x���f�Qdy��ۏ�ܷ�s��@�2����f]�$�gl���t(>��`*n��r��!~8W�������s�T_jv#/[�@�isn�1>��8�*�����?@�PgR���]�Ӽ���rg�8/�1wy��u����̬g/��t&A��D2'���+���?�x���b�F��p�-�i�/�Z�fK��#�Mدlz{A�����;����k{r�,4�U��^�i��?O��G�����"�k+�(ޚ��:�m�9�:��W�uH>���,����݉��Y�J+�a/�*C���k�6�v��n���������]��^�%rY/�����Z�L��3�5��<�x$���8��z�9�ʼW�e��3 J�ڛ�V՘����3<�\(�5���,�6�H[	��\q^y�pY*����$@p)jml!�JTQ|~��ަy��<67m�W��iN��.��JY�@x�����-�?�����OᨡQ����0=�@p2����w1��7R�������8����-v�7��ʅ8�O�Ȧu�=���a���A*�ס�MG�E �L�m��V��,��j���ƒ/s����T-��͏��x�y�j)���2���^����%+|�W����@�v�B��6!3�!�U���,Fi��)���7u�٤]ʻ� r%"�����Nd=�0���J��kZZ���&v+k|�+7,\���RD����љ��0�m)�b$?V��������L=]i�7�j�X=w?o7F$��x�U�eTbǕiKE��Ґc-Fzk��+�N��uR�������5��p�m�72'�r$�W�XOʦ�Z�����+0�N�&��ۡܝ�)�R�f�w��3{FZ�����֕ɼ*A�"?���i	�m%��ȑ����0y��Yq�9ލX����͆Ô
|��s&��:��]˭""��c�m����F��H��z��Bぃ�����R�
�ي��.?�V�[���F�)y��*�����
�՘\�pݪ��-��dXYm�dO\�bUŷ���W4s���"1CW�#���a����Q�O,��\+(�x�""����󐅰���&3f�_�)D,L�[a?���PU1�����C�rzH}!������Q�
��o؂	 ��e�oH�0}�5{���S�]b��:PD}8�y��Y�qL�Klo��I.��j\�t�ȯ7�G��1)*�~d`;�5!��'���T�d&�U{Dኼ�7{¼G�!�ԫ�����w��N��o���u��\D�d��R�⣎�|���jq�+Ĵ̓��s���t�RN%r>��:3��a��o=u;X�%�·HYb��j����[V]��|b�؅��C���5EӴ�*Kc6�zg0����~�p�G�2��*�j~9�²ﵘ�)�,���b)υ�<����S���m
��I�ǶJ["�J��~����Jy���f��fӌO���)�zHeZ�wUߟ��E�#^I�:���c������0��O�O�gu�,q�`J���X�	:�7l���7���"�GߜR|��<�����o~����ŀ�Q\`�8��A�0�`:̞Еvݙ)g"�޺��0j���W����f�g���/��(J���\�@=�e�K��Jo�0u���R�[��w �yn���E��W�<��󄄨��V6P2�������Dk������,�S�?���f�H+ڑ%P�SM�j���j�q?|P��U�:�O�(8�˫#�8�6�/켌�\=> 	$ڇ��.�G����)HJJR�s�j_lQR�98�#�M���\�22�� ���<��UUO	���gQ�I!�}h���{!]���@�Ö�R���0}�K�������+W��m�� �&+���+A��s�;c�����id|�\uļ�E|x���I��-�z��\e���E�_�05�����ݛ��rAim̄�����C(;������+�G+�xv��u$�8�,�N��-X)��x�W��x	oo�w�����@nL�&z¥���uj/��_�7@xי���s�H��l�%��� ]���S�v��>�����Z���EAB{����:�5��v�ih���
x�~�J�i:����%~��x�Y�	&��	�~^��2!��5�_7���Bj��ȓ��]�'{D����y;�. �rGnhُfln�[���5X7���kI��N�]*�V I�p[e����Q��A����/>�߽Z���=��
��Q=M;�?�����qQ5M۠"(�J%�H�9����3���d$�#�P2�$I"9�$�"90�9��9��~O���w��ﷻ���8�tw]UuUwu5�;q�[|6�)[�7�!���ha2�V��1_k�w/1�Έ�)f��))п���c٧�@B9z�;�c�D-�g97~+�wo�i����ЍAo�Wp{%a^c.��r�GV�
'�L�17[�N�^�0�~��EO�6��^Ͻ�x�=.�C: 8ͭ;y�L�{�쨒by��DSya�B�$T����*�h�10o�(:��`�K����h�P�)�7�W��p_�;�z8^�>�$���}:Xp����X�XpQ�ߴ���H~��Rnt���:Y��8�g��5T
n�AV"s0IV<�ӳŲ����������9t��o?�!��F�$�~�FU2��'���k�0<�E'E\�=u��.#��\��];ꄄ�f�=��x�B|P�dGY���fY[[�HOO����z�iڥ���j��His(���I^EFq|�HY�3��ɋ��ee��ͫ�fp��gΤVV�$��[��X����  �K�W�{��vW�:��Ν?/���+��T�����6i�]�P���.�ф K��`xx�$�2���tj�HZnɏE�x(���e$�]�x�ů]�$E|���.��˗/�WS,�~x�d��(�1�*��]s�'���R�p�m;�#�M��"� `��+%%�{�b́;)n0N�++�h4����ϖ�N��`v��%�0�N>�]��44���}�+�b���cڎph�L`�K�u�n ��/ǃH!�XxEE/����ND�0":;;}y��3�lf����w�;��������EW���gl�>�L�����}K@�*/��§�����!899����yzzJ3�t��� }@l�K,!���À�H�
���dd�0� �R�An��[Ź��
P}�9*��p3y!/�X$3zN2(��L �_Xh=S���5`�oĭ˿���
7��P�O]Ӂ=�Um=�)��M��.� J����`�߄)��ڵ�M+�C�@�����7��u=���ؘ�����^ZY�L
H��QbWJ.(ࣦ�f7Wb�>%4��Us��2?x���s�1���U���
���j�������ɵ��6��W7/>���[��f�-D`C+VV8��L- ��顱��Z5��y�F���[��k!���/������T�_�����KH����x{{�]楣�{]t�:/
�J��'�OΥ��K�� �}�����Z ݇��q��+߽�
����~Ր^J)É�Z��i?��G�����^Ⱥcjj�5�Q�G�V���=vopÓ��6�22�tw�]d.���m�׊���Ԍw���+Y�6����6S*
��Ћ@�{h�|���6eY�E��p��=�t�j���E��yJ<�*i����B�3m�W�������H�����=Je���|���3����E����n:�ڈCy�+�L�Y^SSSJa��.~�}V��� e{�6CYɹH�y>;;�UO3N�@�|Kn%�W�kz/��$`� ���Y��ӊ���������9���&�����w&DgSE=j����OM{����~��.j�s��Y�Ą����<�dж�����rGR��B�Z����`ֻ�]��֖^��;FeE7G�dޭ"����*X�jCs��Vb�}���(��G�ᗑk)�#a�D�K�Ї����]Dˢ��mO��!�2h�_�����~�عv䂂BCC}]���6|�Iy}౱��66-���
f�7���P���&�~	'(i�uH��.0l��u��r��]y���
��f��}zVPXp�̧��<���V�4<պ
�Vj%�)��v�aQC�V=��ߝR��O��s@l/SG�u��u�J���'y���/��\�/f�e�7��7�k�t6������[!AzԀДQ�`�gf]Z��n��_��9����n��������EÁ��N�^�"�B�`��u���'�����؃��E����> ������)�������������� ��'���j�b2nTw0vM{�[b��N/�4����ù���:ӑ��\g�L�Mfx�%6{<7��$�q"��F|��*�J����%��~���P��� �x����a��Dn�&�9�Lː-���OeM�${����T�Y!B&	�EV�\Il.�v����N���ľ��z^h�Þ��97�]��D��UW0Kr0ʐ������~���j���Z�{ \���(@1OAA�:	�\!!!�4��"nO���b�����dve�
0�<�q�!40�<l�L���u��2<�� �j���
�v�	G���h�N��O�Ү��Bz�_�G����W|詝��p�t�S�NCp*�q������ۅcaa�[�t�yWj811���[�r#�D]!��8�g������
٭%)^T	����"z��v�Q-���\yD"H <�U%9��5����ߟ��6N90�:����/�+���;��Pv�ݬx&Q�r��X�｢�6#4x�*�'zFF�d*+*n��)ڱ�47��^��@��"�ǯl��ͷ��Ѭ�Dj����������͞N�Zj)��3iĻ�1�h������(���5]���#=g�1e�ؖ��$Uϋ�*1c5�k=d^�p��oD$�X-y����̯�7?���BW�[���c��' ���焊K�yc��D	�7��W�]i.�E���:���Yq��a��C97���2V�Vȷ3�b=<�����v�4����x�~�]�|���#( z�Z6QF8U�\]��!�]b�)��m�++��"5�b75㨑i�2,i ���{[�B`PNlmk;Lq��H�y�ϼC�;{�(Ƭ~ǆT����q�A�����	uc(����e�:��W4���[2r�۰��R^�����4���
��^��j�ܵՖ$�/��]�2�
�s�M����Ö}���u�W��$:YG6����Ea�(G�ޣ[w6W�m�}9kܶ��Za�������x�G��_f\���K���7Rw����/�R� pV~�H�_� D�̍�j
NEES���i�a�|Ģ�c�;8~�5�iV9���R�l�ֆ���8OsL囮�Sn�h	��G�F����.P_�{�T��v���~=˫dn�+}?f���K����e~� �ݮ����d�wt5��ۆQuQ�P�g-�]�qon����c����
ij�=D{�o���w<��^Y'R��Q�=�3�gBF��bz�I����ʕ�B�Mד��,���}�VX৬��j.��r��!�:��'d#`_��@��ȕ�u�>yD�q������.mc:a��ǒ���VaA�P}��n���W����ss� ���$����ȚnkZBƨ������S������sG#6��@�/�&��n�p&)�2�*{iA��X��GJJ
}�
�=8���#���
����B��3<\�qѲ��]��}zA�3�AYU��`%��|YҢp�&���E����I0� �$ݣ�"���mO#��b��jRXFE�A�ݜcŰZ1u�c�W�^�.����T���w�*���0������nV��˲f&�6(a�"8�����f�r۴�J!�	��=�УlyS1�tA����="�mh�M'>�W�Qo�ӿ��'�~����{��}������`�I��Կ��F
�ኟ�@�V�$�8�,M����,�����,��L�ڐ�"�X꿙�3�gl��%Ľy,:���ꯆ�!!�ݡ��� "bΏ˼������j��IX�^�`w���)���H=��	�	��E�^�n#��+���h+t�OY�,�_K�Oury6y��Lt3�B>DV�[�8V0Sg�[b?�w��X�.H���R�W�%A)-�H:����~K@D <v�}�C����ksW`����0�S$:3�9�B[����ٮ�D�{*����}P-�,��Q��ʯ��D��0�mع�+�9Ϗg��H�fc��lmI:`(̰�[U�c�����i�"�Gg�غ��mAR#;gf�-��H��� ?�L���
����u�E}�@/٩�S��R�e�}��Q�M�,��3k�R|���O ���lݹ�{̧�����ox:>��o���iWJ���	w����yq����p>aa�Y7ps)}d'�x0��e��Ql��ˀ��|��2��q��uC��^����O4V��b�@�>��3��@̼�@?$��������X	0?b_;[G��x��=��i���(n���{;>����T~6�`ફ��QFw��r�-����d�{�a�cQ���rི@<�@�Xx�,bZ�55�,1x�&�����qh6#9��z1� xβ#V赤'��A�׻�qP��XO��ŕ��@PhYޢ{�u��P�T�&�!$�3����?�IOD�~Ry��Wh���Q��,�F�yhN{�������f�e&P�q�9_3KK�7��ܘߥb�byY��;:::\cG�B�o��P�j��g��0ν1��9��W��%���m��QO�F�]<��,^l�e��p�3����;���)��nqwa��[\\��4�Gy kW��(�)���u�N{uY��8�yv�pKHF��PoY );������ĈFĴ�ZEyy��;�<wd�B 4Y}�ށRʈ��Vo�;��[�i��#y@(.��gt)0�h�wV]V��@?��o��_vF�@�{���m��Π��7o��\(4Y�V��"���x���Y���aj����C)G��?�3�<�-7F��
�q���T�j}<F0u6ǰ���g���؍D����%@��]�̀� h�yg�7B0'B�T�m�"ȟP16& �������`��%ß�����QDu���KGVUx=�LUN�9L�F����v��Q�75���܇��G�~A��L]����A^8��3�V�`���!�������[�����Z%����^���Du�ݳ@ ӌnf`�F°ᑯ�2R�Ү1`�/�8��՟��#*G���:�)|���ZeC� ��=�����ɛ�"�,_�h�E�T.t$��Z���{ݺ$�����x�Dn���f3ݗ�/p�`�b�R&���b!�s+�"�}�y�c,���	
��W��3t������qȗ,I�'^ 1#��@��EL{�� �HT�g"�``�	;���@�6�����Z��BV����`�a	�ec�k�4�#V D���w�ǼP��YJTz���L?�T8�d�(?^�ě�j���qi�����H�9A[Bo&6� ���%9�c�T��r��x4����=�"������?1���Љ	�n�_��L�'�r`��u/%�H��$n���].��B$Y��F=�|70tN��"�W`ޅ�A>��;��X�y����[��	����KNe_�L���Rz�U�7��lB��d 3������X ��xW�gX&^�e|���guk�]�y^��{)�©ǥ��X�o�f��o̯��ɧ{����|LWL�J.-)q���y�{�@唋��@� ��3�A�jia��=Z�����aEww�Ej��_��|���Li�ۦ�P(d)���M �ں�u��r��[v�/Z������^f4y����Ho4��K樘�
�w�n2��n�M�+L��bRrK�RU˓�F�� M<�:�sG�?gmu��r|�2�Q	��o�0Ǟ�+bt��\�ỶJ��]k�ύ�5<�F-�D�M��E��+���1+q��;3ƇE��� {8�{���a���~��Zz� ���~��ӿ7�8�~�F:�1��]ч9bhu���x_�ǜcV��ǆ+|R�}3P�%?77���$vy�T��jտ�7*w���j��U�3�<�����\i�!�)tjd�+�)�=��4+�G�	<��d�f�̢)����f��U��X̪���1{d�g�m�}��dI�n��鳁�]d2���{�>���1�z~x��QE���n��]�O�4����g�7��Fy�k\������v�ü��Ύ755ٍc�J���&�ϓ�^烠S_�,��C��SFRw�����L���uCz�J��˧Ó��=1�����;����^p�9Ǩ�?j�'�{���[�zìC
��]�*	�o	AW����܊�|�����\;���ӱ�$ױ\r�@�n����.�n�N!V?ޯw��M���@/Y������vq�|���r�o��)Z��h���U�+��Q�y�+�mQ�+N>#���++�AC��B��n���d#�ܫ^DwYwF=��j�Z�����؞
�������������y��qUL3���o�?����sȾ�i�cƥ{d���^���Sl��n���s
vV˂w�����Ƚ�oyBg��u~���fT$��ؗ�(~m��xj���L��<G�v0U_��ͩB3?��(?�ۙ�B�"�͛7{{{�zJ�a&���i��%��ٳ+Vl�W�0�=jt0��TVnS�ٙz�4�F�¸$�gʜr<�~�1��L���.sN}ɲ�'�������a�n�a��]�S��0�J��ג;���Q���n��-��]����ݩf����μ�85Mj^7�[�WiL"�##>�߿� ��� W<=9￞?:
���N��B$�M��V��A"�[����t���O�+}�h�������w3r���P��}�����+k�q|��fgga��vo]��6!�\��宋�&�i6H��Te����c��o%�Ku�>�H8g�شvc񵢕�xQ&FQ�ݝʘ�y	��,�uM�����wFJ~�H>��m�MPH(rC���0K���/Ow0Os���L�kũ{B�����8;t�Vɵ;of�I
m0�U,k��%_��L��0�so��8	�t��>e������/��V'�p�d��-�����=�L-8xC�ESs��G0�u>�yeӽ����<"�[�����?]��H�k�9�>V�.�����)�����0B��˗��\���<x�}�/t�F���
�G"1I���ͅxIE��k9��>�Q{��@�.����s+lg��@�I�3�gɩ���/d�u�b��>���/&���q&3\�9�8o;\X�k�E�А����Z5����h�;NN�?���o�uw$b,��EP�����7a�Ű��ߏ,]�m�M��C]�]���j3$x�u��$���`J��A4W1�΁�H���ە�Ͼ뙷���E���4455�*;,�;;;yTȽ�}��|׹l���yU|����0�B�`*ƴ]9M!_Z�S��_�f�LHO����+���Ƅ��V���+�y��h��s�1߆�C�n�'''	]ʍlk�Ɂ�L9�Op>?_�+��UV9x��Y���)�.t��&�`�!�b���]�RTs�������	��8����c����ᕖ����gf�310�G�X6y~�����=����:���eG��JϜ/���J�8��sK�X�z��C�|���5?m�3��Nt��~��=�H�f�c>\�]���4�)�s��c��V1x-��� p��+,�=Ӵ�I�x�ϑ,���v�d��Kv����$��_o����{~�!���@~�Į�`5���L���A[*�'K �(��K��;8s.埉f��;ք
��}҇a6�K���x�&ċ�����Ψ �}_��W ���U*�y�`8�޼@r�)���J�q�y��_����.����7����l���i�f���e���3�b6֮S1�g���޿�2��_yS쵍K�o�q�u���#��{Is6�0�IArh��'+I��-�i�l	��54Pߞ�r��{���ݰ�����g�w/�|+���	�Eccc�M����L3x #�����؁ϑ��4=Fc�pI9�Xr���=!��e��{�~�̶}R�/�o?�߷������~�O�gS�8O�F��UO��=�_:�����������CTQW���僱]�Ī�4B�?hHYh���5'''A��~'������w�3~��Vi�g�z����b�i�]���ո��t"�;�PhHȌK�Z^Wbq�Ư�]���7QG�(�Ra
���W8Xg�ð���;�4�$�67���*�I�(�����H<���|�۷oo����&Y��L�i��5�=~U�B��/����bBT�Z�1*��u1YYl����AvVn�=R_�6�f�>��t~i)��K�}9�9��ȍ��T�G2��{�ĕ:���Y���Z=��U�d����#�p�EZ�v�G��i��m�.ķ1�!CBB:�vV��y�f�W�9��W�|�IP�$��^92ڂ}B9�v�?w���y��.��A3��t�G��.�#w��gm�����&�ĩ��J��%�hٌ|L:��}g7ջ��"0��9���[	x��y.#u�ܗ��)��\�3���:$e6[жW�?ǲp�~���0�={�C��0kX�Cs�)և�}`:|�uN&\�y�<A�R-|ܓ$�c�1������O"�-+2�+!�>'���9�9OkE"�ͣdIR%����� �SiuB���6�(D�3]Fܺ��^��R��a�j�%Ϸ��p�v���n�t�u���٥n��:��nk4��@������o}u��Zʹ#�-u#�g���f��Ƒ�l��;x/QOkb��� ��l��<5�gѓ�*թ�6��| ��� t���/4`�:�3��kt�٥Y�#xR��6_/�O�ʓ�Q�1G_}����ma�-�9��\�˨��*T5�������{�͍~��?5�z��"�;�춨?#_db�z'	���1u��	�!���Yv@�:�19Ɵ�D��-��֤\���H�҇"]h�
���4��O���(�`M�_�e| �S�^��(����0X�(�ڭ��d}��U�驘��'��T��8͡Ƶ�_H�3_ν�R�4s��V\�mAfA��^NO
���P�"Ab�_H�����5Ar�^6����k���]����¸nN��?�e�8��#������NC�� ׌����T!�R���}��K�d�˶c�� ��>�s�	��9I��9���.v䚜����_��)u�s�0��ԟ?���<Ir3�Q���^awg:"���	[9P�Q��Ŷ�6뫖�������� ��� !��a�8���
�|�T����uT��L�^��:��ź^�tfn���؆2F(x�w��KK���?����RkW�7t�z_�ӛhRg�Yl�G��$��J�h+�E����\p�*�y�|�Y�5n����uHT6�x�/��Gc�_��O�=����(`�2�~`I��V-hc[ڤ�ov�?d^�2=m��+P�H��:�n�׽p~_��^ ��ζc������N"�<�H>�~0k|b�h��c�zG���UÇO���D�C���1�X�������V��Ns7�v$�����ǥd�9�@c	���v>
����QMJ[#,**m�������:��v�R=6�Sm�n�9���Zz���D~��v�$�qt�#�����ڑ�P�U�1��M�����~�tL��G ��/��-��L��4��F买�i���j^9�����ԫ�s��&�J-�ЂR%D����6މ�R6B��c��?x�ݜR�����5�<�`]��gR�P���������޴>��B�����÷S抭�B䛳9NFH�5t�5��S�Q��pc&r��)7l|8:M*o7�seu'�t�}��_6�p�c�~G�\^R����f������ƒ*�prY;�2���"�#u�،�W4��%:^���d�(�ɱ��wdS�U�V '����<�Uf;�]�<�tS~�~���E�4K��o�p��f����&:PH��U� DJ���X���+��0���*z��E����7?[#o��%z�ymq]'ʮ��]���v�Q�9��	�-�W�tj���j)��DE:w.�5��K��������a�l=G��r�ށX���Q�`?79�9<l���wm8Q7j-v������퇋ٸ��?�d'hHM������E���7�b��N��10sy����G�X�M���*�iP�XV�l�.��Y)��j�mJq)qq�vWN⤑|_�.����7��>XID����.�7F2T�w&��ǋ�64�; �����Z�l��y�-�j�:Ue�+�V�Иa/�w@57G' i�}���N�(�j�*!L�[zU!��+/5���:
l4'�#ߴ��r�Lf��
 7p(cl�p��""4��*��<sD`�g-݈A�2vޖ[�8ࠍ��!�}y%Ɛ��"s��wV'@Q�5g�l�(x��ۂ?��¿

9��{�-��m@��s�P�Ҕ߭��j�5`u�R�z��[�l�׷��9#xpp[Y>��W��vϲ~��q�	z%w��'G��V�i��qД�ز�i��'75�q���r��7�Q�	e������+�Ȫ���<wtvK�įK�^q&�Q��z|A�2�Y]�Xl�?�F��$�B�W�Q?����`-��ￌ�d��Z~�/|ZWv���95,���M����|��`��vwy;����J�ƭ���}Z����s+/h��nҊ|Yy��������&�<݀��W����V��5��Y6�7'Qd0�x����uQ�K�r����X��ͺ2������HT�Tqpjnjn�&�1�
n@a��J���#�%�������ŷ1̀l�_G}�RH~[s9�C��,���l��jr�����O
Y(�1lOd�b�h?mݍ �;u`�U�-��{�Id�MD���Lv5n�`���1�Yy��%g}�Zܧ�|�}W7x��I���.&ҼC�R��M�w���^�>���[yt��ݑQsIbk�u(���Cp%
���fT�#���h$Ms�T�ݰ���:���~h�$v�;�~�~�`d��慝�`L�;U�3��|���Z�l���η%9].���U�'�lϜP}E)f��]ۧ �_�<Q�����>��1�&^$�!/�[uq���(	jJBח%/�Y�h?���r�C6�q,�>�We>�c�0�����ӥT�ܾ~}r����s�U�卉E����
G?�UD[�r�a]%Μ�����U����Q�6��b���Zb݃� ����1���c ����&�yN�_�n�]P��7?���nI�5�]�˲%�9/�߰���T�ϳu����x�J�gS���9@�eCΪ��r���wYܯ�"M X,ԸG�h��3;X� X"X�$����[���|���un�`��}I������a�P�oϚI~)$>S+d�nq�7 �������mh��6���,P��uam���y]c!�.�>�E!"�ɭT$�Ϊ��0`�Q�Y��0�<K�u�X�Z!�mAʢ&&H&2䵨\q2�7q*Hb�M����&�yw7�0��L,��7���evz���{(CT�3��)d���*˓@U\��~X���b	����D3��$ !�x�wv�Et��=F��Qt�Y@ Ae�qO�c��_(P�v��F�{m`�ԏr�^H�qw7������i�����B����x�=P�ʏe;�r2e�A#��RH��q)t���li?���дE$��[ZM��QɞW��g�h�·Zʃ��}pP�w5�:��48Y�lZ��h|՛ cع�.�����)i���a�M��'WQFqްm�J�Y'G{��X��y���4M�	Gh�_(�'İ�Ъ�|��o����Ν^Tz�:0��5���;0J�jlΚ��;�������!�w�O3�g�����ht1���b������$UR�>�7:1h��3�m�9���Fu�f\H�Y�{�RM�$=��;�,/5~����)^U��|��3��R�+�~��(t4n�/��d*_:��7����΍�� �LŊB�a' �tz!G�Qnh�����f����ȫ�c��#z.�.��|=F�(0jU�3JC���Ű.	��k=�����������W�5N��g��.<V_��u)�i}�k�'֤����Ǆ��po[�2Yh  "@��K�퍯CC�?���=$#�z-;��A9"H/Euj��L�BcY��;�.�9�E��9��Ft�A+F�Y1)�@E��d��_�&�,�����x`��e<b�����S¼�œ��ۏemp=V��FJ�0�\��m�}�lM]��U�#�f��F#/����b��fOޣ=zM8R��3�>(�{�V���GX�
�������T?���C�4�&����p�c�P|I��@���5�����'\�9�u��H���עQ�̸��M�T�i��S���|�x��tM��Λt�n����v3�esV�@8/�)�h�5S�d���M˄`��>��y:��PI����]ךz��/~����vm.H�ߛ7�.�u'���1G<R'�)�AE��W�$��U�-����)�B&�X|Di!Oa��H�I�JE	hKԛU��h���Z�kNRe��`��Z�$W�zq����\���m�'���ؖ2��S��[A���&*�ӑ.B��9���H. PW�߿4�QJ
�F�3;x��˼���eU�@������U{ɀX��X����ɛ���u���$Ͷ[�V~��7XQ*T��l�T� �Z'<�#�2��.5b�'�;|�N�ȼ3Y���j
�f��X�r~�@��3���2��d4M��:�����=��~���?�?FE��BJ'��'g�<ēuq��jt��!<�c6H����T����'u�FP�}H���q�
P�SN�
>sC	�{M�c ْ�e��T_Y-':������&�۶%-G��'��O���m6��fX��;{8�zs�����G;h����=44�|�o��<ړg\i��6���9Q`��T�2��|/_���,��q�5�krӽDԐUҲ�sD *LF:]=��%��0��PP��w��:'>X��aۧi�}4�/��S'q� ��9��*��.%�&�\���.߂�Ǯ�b�!���S���6��g���P��hI.z�ˮ������9���L+��5�f*m���xIu����?f��3���}_2��L�3�2jH�KJJ��Rjv� wo�\���^�}*����fҞV{�X�H[�5����F��@id���F�{� �I��T'"�]ʽv&�[�U�;=�n�DhdC}�h�$���ۡD����Q�4o]��4�M㻴���+{�0���K�];Uf�d,WL�`T�R�З-����n�іLװi�	�	�����^yi�UV�$�sE6Y��M���H�'������@�{���s`L�c��Ts0>	�6�Ph
b52�A�����=��H�1n�ݥ�����m"����u��q߻�J?K~��/+����-�VK;zO�V{z��P9nE�h��(��֏�G�s�CHq	���	!f(�2 �o��V.T�Dg��iYi�%NH�<�٨��Qew�7c�d�l��fj[%��4��;]�C0�۩����K����r��jߠ�Q�¹�����4���f�$��%KB��^��Ɋnp��T�Ǡ�����}���W+ 䉾��Q��1��K<�6�=K� �7hA���K��}����˅S+V���+%��G���7\� ����J��I�/�����[��:@h�p�h�U����j�L�J3N�� �$N��=�}?���̖)O ��߁�z3�%��gj�~��l.d\�f��ү_�����P4�h�ڝ:^R��z����U���(��0m{�` "���M�3��`�.�b�P���zm��K��W�j,��e1Q�G�+�A�]?{��m�ڃ�k��u-��ۜ*��)&-p���೐����$�ܰ�,�j�C}#25�V88pM
K���ٸ�?�#;V�hU:~6ǴV:�k*p�\S3p|8���e �W��8{[� �$_��}͓}��E psp!ʾ�t�Ͳ<��R>����z���o��w�Q�-������U�Ş"����#��ܴ-���kz�@��&>�8�	$�֎y9��ok������h�� _W��+*)����)/����[����J��Tȵ���-�����k>>����%~�ZA3u��.H���u�~������[���㉭��ռ�u�q�����Jaz��I����6���L1k.��6�^-���(�?b2�ߝ99����<���E�c��9�?2�5$���x������/� ��z��iT��О$#3�rU:cy�%�N{�>Ѡ���j����z�.3��m�B�\%�*��m�bqMS���)r �L��!�4�YX Y�I���`IO���sK�f�@��۔_Y���ާttt�S�;��`t����1����N���o	�+��ST\��%�.�yr���m�ۃ�ɳKx,}����,q0�1��=XC�:��fk�C1c ��׭�����z�Ay��������\�D��6��A��v4Ĵ��ڶ�+I��q!
~�+�X������ڙ,Y?�B�Do8��-���`�
�P�YD�@�,d�W̪���c6 /6.�b��ӂ{����BW3���ϻ)�V�[�� �\r�42�<��:=)tx��2@U�ƞ�B�Db�� ��	a-�p7����k@RX�Wc��6�v�i��s���ɫ�B8����̘���-��lj8�!�Sq܅��!���H�pi��A����a��\�C4�����Ų�X���!����I~���O"Gǃ �<�{�钾��n�Qr0������~[��up�S՝I�H�p���ng���Ǭ1P�@¢���d�h|ۂr9��7�� :`_d����YC�9W�hS�S����R�	r#���ec�tftG�J{�������w�A��F��0YVU$���0�R�뱵+r�?<$��¢�i��=%��i#�[B(�Chh�Y� ѽ&	�s�`2"�B&�+z'�� ;�&`�m[���K
�+-6(�r� ~+(��
:�*1��@#�U�ǲ|�N�����p�� �����J+a��E��9oe��
M~�z��'#q��/i"E���Zc&�i�if8?�C3�� ��?�F{<5֟oM��;ަ�|�GA=L��������z��Lk��$��Sph�Dr@S9�gC�E1*��n;K�Gh������Z,��Q� 3�Y�������>.�?	)rv�)MKw{���BZ*�6����ii�J��VJF�	��[#[|vԵCʹ�&Zko�7Qo���z��ik����%R��M~���Z�u�ߦ���(�n_NțƱx¶K/����M#���&	<�E�����9�J��+�7���&Jj���Z ���n���nB���1�q��qu����rW+$�n���i:"N��d�ZA~�K�-�0��J0M=�63E�4ޕV�xa�b~��õȴ�
d�� �FZ������Y��ЌnK���^/J���S��Ē�\���v����&U��^�\?qП6f��PT����_L���,$�p\�D/���q������Y�^�鿈��\�t��S����9BG���]:�b�M"ty�?��B�J�v�mi�
��.R3W=�}��rN��5����^Y*�j���h
@67��)�~�q=�%"%(�������0���2S���w�iL!z�#�+w�������R�����}�Y��j�f_6����Xg��j z�F�������?!~P9��/t(�_����;PI��o�q�K���(Wsk*-�ݢ���]����R���@�FB��>r�>�z@'�cp�HKGB���d<��l��i�J.)$�f��%	vP�?���A��5Z�xMO^���4��N�LWY�__g�l����qZ�'��W/'#n�NS��k���K��d_�ybNz�?t��EWVC��p ¼�?���?���?���?����g@���N큚�D�bm�H i���l1�����>�P��m%%�}�
�~ n���t�Պog�FH��9���Zq�u�Y�L��L����z�6)1��	���iRX����1��J�z���E�����~�\�ľ�dF��Q��K�jvKɉ�]��j��~�Xt����=����h�Ց���:F/f�-+�ܾ�k�me��h.�%&&x�-�BS:E#�j���do�)������M3�?�f��~�	�"&1a9�`���su!�n8�Ӄ�@��@��@��@��@��@��@��@��@��@��@��@��@��@���CA)k�C�2�`��S�q;�g�!�?���m����:Pb*wG
�;��H���-Mc���mZ5����e�^O�ݗ��8����]Y��P��5��֛-��	���;}�(2�sϓ��Aə���6��2m^�Hb��]�Bқ��o�J�t����A&!!!�;��Qi�ȓG��^�'e��\�#���X<��|��o���^ �l�2��ԅ��SP��=R���#2�ۺ��6	�&nyv�md��t��9l�e���&�r�����<�r�[p��Nv��a�_��FV�-w� ���C(��p��|ˣ��+��_�ݴ���������S����$�]�����3�v�n�@(K�_�p��Y�լ[4�Rw@���>T�}/Kr�u��k�j�[�����U���,�,H�5i�1t}9B�z,Tj5��WXg}�|sJP�sS#����>bA�4<8g�Yg���:�K��g+D"_����aǎc�q�q�֖����\F�P���S�
��9�e�ڪ����m��9��'�H�Bw�dV
^ ����s�l܇�+�P�R�ݤl���ѹ+�Ji.m'bL���YE����p��b�l�h�]&�o�W�!���'#���VRÇ[�mU,�Sz}*��ï�i�J�k�{p�Μ.�m�����ݢ$��Na"�́O��?N�3i��d�q�׌,{\�(p6tht�eBBBu�(z�q�\�pG�\^�9q��	ua�	G�Ոj�s��Z(��}�u��B���n��fkn�׿� l�����o���~���h�z�FTzw"�;Sd|}<@�OF��qx������p���_�|%����@�w��ǸJ�G
���rf�?[ 
Ed��t�WD4��U���yɻ8c�"�����m��UY[�i�DB���K=��5�?�l��o$}��G��q�ޫoq�Z8n�z���fr8���vkw�����۫j\���guj)��R�C�F��&�!�4�
Ѣ���_����5rjྫ*ؔ/���)�M��H4�gO�~X��Y!.,�:����c��4�$_[[���Ms�6��=T�	�n�y�Ǖ�����8�t��s�l��×�^r;Ǔ ��� �O=P5˨%��oE�.����4��25���/8;���|&Z梵CV�ߵ ��|��U�}����mB�F��>������m�zl��6Ҡ
�e�m3p�V���א�-�x���ZG���]-��Ȝ�Z	�R�(Ԅ*K���`q�T���sͻX��z!Ii׍/��,�^�ʹ�Mo)�ާK��]�A�[>9/�:n����T�J��J1J2���F.V~�2����`ۣ������$U2S�����i��Q�S�����x��*�^j-t��t���	�{������`�Ō��[�}���������l�KK��� |TP1�����L�j�햋E���7��OU�͸-��N~����'�6T��B쑭E�b�~Փ\4(��h7��ܟP%���`�_���y &�����Y]g�ɹu�6r��cL�I���)�=�����u�9�.�9.j�����c�fi�C�y�BB�Z��}P]Æ	�"�/��7�/���-n�� x
ru�z)��O��o�$�S�R,�#NXZ��B�9��6�����b{_GEYC�pF!"ۧ�IW��p�s�r)�&�L�s�3nE)\�6�m��@�s��!�O��c�.«WK*�p�I97:�=s��~�'����<��+�z�_�_c�f1e�>�n�S��uf�GG9��\�W�@4�fQ��F<`����e-En�WK�/��L��>T{���ث����������#� H��A�R�+��TCo	��"]�w�J��I�5@��B-���N�;3��3W�y/���s�^{������Y��F[Nz��D��|�b69C���G%�zz]�cu��R򓍼�x�k�~���h��`�yѦ٦qp}���^�j{�q���������缧dՑq���w�?�P��T���\�9� l���|5f�̡���7� 1���(�ԟ�����[Gmw��j.������@dZ�MѼ 1�����0JA�����j��T3c֐a�Y`g�g�o\�����Yz�5,�Y#ACu���E	E������QS��]��h|�s�Ƿ��TtX��]��X�՞(�?��z�L&�`G����o{��>�g��D� f$�>��s� 8�ܰ �S=A�J$���6x��q[2�U�1�Ñ��ٸff�V�XY�bW:�M�d42��͉�8��=ؿq����}mm���Qw�Ӌ����;�o��P��董o��?Zb�6^��M7��J<�.��d0m0���d,�}R��Ҙ�g�Ѽ��\X�(�횢�#.�G�uaC%���rc"ڼ�0~�t;:��'����\�^Ɨ	�؄���̉���f���H�U��Ő(��w�N�;��V${�y��c��ۓ�����tJ���8��No�_}c���r��|o�E�����eiQn���k�@L{x4�֭))t�?���u�j8���S9G��@xH��5rz��[���#|n���� &�s�M�o���;��:P���~��Z�O�4J�#��8��9� sl�YA��wNRE����kd�G�R\��U���b�a�>(]���upyvt.wH�s��)��"@��fNSΗ�)��O"���o yc�o�yjg� ��,����l��b�D�O�S|d�<�&�W:E`�~?�v�J���1��d]%�^�4;�ͻ��Uꏇ@dF�5S�>���ט�=$��\�i��)�D�L�	�By�¾�� ؃m��S4�-r �C���ClOR*�s���=C)���]jϘ(�<�����r���\Qq�Xx�n\�������G�����4Q���t�T7Z����b��&��֖sq{$9�	�����A�!��hرɜ$A]�{�2g0���5���0*CR��7����Ӗ�tzڨI�5۸~��q��T���9r�&���d~�������7�~@^���Ɖa7z��Yh�Q��j8�A�P��*x���EB�`���;�Z؏�Z�)ۄ��s�s�(OK�˟��D֣��_�gى5f����sF��Q�Y�����g^d�:|����:�>^��R����½[l����&\��3�h��SV߉P���IK��7R�)}s-}5>e�Qfڑ��X�`���X�$�V]m���V��C��o��.�%�fa�_�|�����gO1�'�H:y�K���ݢ8��;�ʦ�2T���b��q�)��'��Q��͜ɍ?_?�sY^�>�&���{W�9�.�vQU�V�Ʃ���%��w6&�����e#@��7�e���^8'�ᯢy�����=@��áC��C�����y�g�}����*F�WO�9�@ݝg?GyF�?V��6�'��<1l��p%���-w�m¾L�`zJE籡P�s��-J�m��GO1���K��)�}��Ks�Ic!)!!���ϱ�2%B�).o���>#�.ss�������������A)M{>!��x���ŋ��#e9msm�^�|�q���rCܒ,D65o��U�/j��3K֪�����#����[�K��-}�ZRRҬcK5�\��H��/#�@�k���IlV�e�^��|�m�?����P1���:�lF���	�����f#�_�����!���",B<& X1K�v�q�:D%�H���_c���k���3<rD��;�~�'���Ғț�F16Ω߯�ۤ�ͻc�A�i����ۛ�n=�8ҊV/�CFj�ͭ?���쭼svvvsR�P�`��1	"|N�: ��e��F�ު�,�ݱ���,#cb���"�[��*���DWp�!�6��X��ᰠ�$����	JVWﾹ��O����ܫ�;7��[x'�����:�jg�h����t��{�lwsZbyM�>AUQ?�[P�X3L b��R,x-ūew�077����0��Ȅp*zJ�D�ƀ�>h��z����ק�I�	�n���!S�yb�R:���0h�k�������ODޓ�4��XrY6��\��CG�utn42t�1 �9tKQ'�$DR6�ě)'6�+a��P���|ۨ�!�>Sa�x����ˑ��Ղe�	ߜD����Ľ�l�%*�����7ʬ{�rss�̾\?��rz"<�_/��?���_�,A�����s~Ywm�H�=�@��>��+��4]��*///��#|��C�-��J<��L^b����1u���M�}v{{�	k#x�)@G�{����!�����C�U�w*�a�W"iUz�O��\�0�7m�n-ig���RLKK���3As�8���;"t��c������q�鵵�:5/�>���1۔F}���Q��\ ��J����7�� ��N��~P�%.���C\�H-���@	�a�5D�f咿��X��X�0q�ܼ<��s>�V������I����6�w��0 �oc�Q:���f;�)A�+�x����v�#9�Ҿ~�����XB��`Y굣
�J�P+��P5�i7;���H�a�P<��%�z�cbW��/iqf'^��=sGG��M��\�d�#Eb1Y㲶�n`"m!�O�7�2�L�	��m�T!��%Kb&br��H��7Q��@�yכֿ�s�����/�y����B�*�ڨ�=�=����'a��Uy�FD��!�]�����،-PV9�g�����?���׾����{�OKWg��ɨ��'��oeA��i��q�s\\\怄K��}�>}�O�u� �5��E�$b���ղv&��o� +�0̪%��#�T3/S ��K	]�o��־�k�Q1��?��tB�`���Y�V3�� ���u	��s����|�"vDR�A�.L�;S��e����%i��	��	��mmWD[����)�'��i86�X�L �T\\Ad���0o�ݛ��E�v�0�~�G�T�ײz�T��1խ��Y!�j��	�䛫 �*��M$N~�"9�:n�++
G�l�p�q�%���9��(� ���!��S�n��|r��[��%����I;{��k�kU���]U��7pܞLݚs�89��F��\�{�B�sbE&s��1��6�"彔��o|�C�6R<s���A�)��x�hkS�H���I)Zy�zp��/���(���o/�z�j!R˃ln�#�}i� pa��ip������,���5��4M�Xodm����Xc�������2��J:n����Oì	�$>���H�.�/��~f�<�h�	��yz��W���X�'�U;$�If�/7�$WԮ����D��^�X��35� (�g$�����~���s0������?-a0���Ce����IbCfN�Dą `����V��l�i2��(��P��7�ײ�d��^�Nb
B���o=����'�k-^�.�~� �1���(����/�|�Go?��4f�JJ��_ :��Bt��=Q��h
�.v5��x���i3c�D�gΨ���)]R!jᶪ��.^�����Z�O�Aī���!���#چ��|$vu��E�Jo���ƹ/k[x#���2�W�'�r���g��w&+��l�����7�+�x� j�f�v����F��`n A�r���q��>�5��Z�2it���75�bO��F�`e����m�o�p.H�-���;���it��ӳ苏8�K*��l���=+7'm^DR�<R�Q�r��L2���[�X�5�B��K�����{�T��B :"�2��+R�g�!q�7 �Ti�Y��K��X��o�g�~ϋg	�@f�w��`��/(k)��Ȃ�����-V�K�Ŝp;s���[^��1����?�^�t(�>W�Z�����]��v��,�Liy�'=�"�!��o��J�*��B���3��s�c��܍��*�YTBv-f�i�5��<���P�>����*oL�p���n�!D��>I�Q���u�򏣴n�4���6(u�� �]�����,~ʓ��� X��g=������@l͇݉ą��ݍTo
|Qo+n�+Ԙ��җH�:�}qO� ��� �&���!zΡ$��!�~U��!M�u��0>)�΍X��W	,u����������#oF�[�WR�9���!c
�mwH�B�!�}$}6�~T˕�1�����֊��ģ�4߫�������(ƙ���d3���Α �a_�r�T��_h�gl�d�ˋdY�/��9��,)�v�&k++㤓���i/hp:�W[�`�-c�=�}��l���W�:���]Re������U�)����H�ʁ�������E�� u.Нއ�j��g�{���d�o�4U�;0���M��8��o�~�$�	��"��f��D;&��l����V�ܠO�G:��Wl�|+�"�]湊����]�[��À��d�{}��������]��d�LQ�f)�	O��=V��%���@��C�	V���t)Y\Ta$�n(��D��Y5g�s�ٺ����W�)�xP��&�y���:kL^�ѩܩ�-}x�*��\�y	�5�m�.�O��5���# ����H�A�?�3�P���6�T��<��w�/�����"�0���{��&����M�Eڭ��3;T�auP�аKrl��s��*����5r���� ֭�8��n��`Y�(z���nmF�^ݮ�RNKN�Xs�T�I�C6�=�^ /��0¥7aH���[W��ia#巟א$�[��Ы�u��Jq4<W��+��%����b�z�!F����'��07'�,��+�M�m�|܅DD��&�
���-pk��e����6���l[[���\P@��n��٥B>��A�=?��[�����m�T1��9�yʬ�VϦ�͐��[��&>ֳ�b�GF��_�1[Ku�#�4<����^�s��6��f�?f��Lyrw;���@���X����߂����B������C���W�|�n�vqa	�:tmWV,R�����}1.~�X@�� \rܑU�pRH���}�#3>��.���H�����՚t��/$"f�@��vmMb������C����p���ĉqN������re��\���Jyx�}���+W#>C��N��]Ҏ�mQ�ø�pp�:��������gqL]z|<�R�ᥟK[�m�E�D�+�?����L���C{��?�|����&�Z��DKQ=�1
LY�Cm�xa���J�j��Y��]�O�n�Q�$�Rv����%y�����7���N}A09����k����e�(C��``ttt�~�=��u��7a�Hz#���|��īn�
wxe�Bc��V����%�J���Y�r�G���O��{CS��n?|~��xJD�7�H|����K,z�ﾮ���Y@c�s�]	��(J�����?E���/0�)�Gk������r����Jњ{���a�vRW�s��'�~{]�w8�X�-V�A +&���L���D^�����T%tk윲��u�Y|B|�:G��0h�l��Ǜ}��g�$?�sX���Y�w���٤�R���-�^;QhQ�I�X+]sH���;�%���w?b�]�ىq+�����ᝍ&���<:&&I�ﾾ�=C�������\�ܕ*V�8�����|���M!,%� ������`C�I�9��$Lq�	����ӵf��]������x��_Q�����^ �(��	��z�(tYO2�3Æ�>aA�����{��3U;���%�>�K|�>G����^s��} ̲t��6M�']�LI�w��E��n����m��ce1�Ye�̓��+���9�o�Ա�`u;��r�t��Kǐuj����9�K,��y0^p�IĢ�9�y���{y"�q'|���Z���y�=JѲK�>��٬��@|��=���
7=�\/0�N�PV�"��+�K� ��YA�?���buN��3xd(V��6<�[���;��?˲&���SS��VG=�=�1�1�@/�K��ic��揼Q�Q+0�] ��� p�m�-ƕ�Ǆ�U���|���7(��k�ŅzN���Sz�M�a%����2 N�[t�7�98�5�͏��6��w�#d��S�ĩ��:ӹ?�*V;ه�������&�D�|���U���%P���K���ާƻ3Юj�� O版O5���{�~X�x��2X�D#�2�~��	�vE����tq��T��={o���x0�ڠ�k�5�B?nHoo�5
A���� >ص��%���}x�'�(:e����ڡ�u�-�<:��.{���GmKq��q�)L���T��X��4#b���]�xX[I\�z�
7�k
��z��UF���.�)0�Ps���X� ���.����ڢR"�%���1b�p��<;7�뾅���9\h�kא�V�H���ӗ�ON��#+��s����x�l�AaZ"G�T�`�e�9a!�G��j��J�6�L(�8���/ *��9�yS���2���y�#�vvJ�
�kn�>S`Qn6��7�z�X�)�wq#l���铹T�?P��ag�.��"����襍/��<7���QB�sU�c<�l��	�����'��K��|��aW|ޢE��r�%ko�ç�6�v���b<r}~�`�3��ب1M�᷽)f����z�� 2o��H�b�i�#.@���
�K�~3tu?�5LA�H��Z��R}�&b���$�x�_��ym����C,��GQ��ߦ��
:�Sݸ�J}�������l�=6���0)������I']s�W*��#g�pffwP }��͖M	�w-Y�gm�(�y��E%����aҪ]��,��P�܎y�p�m�����nT��ܚ�|/�)jI� 쎍�'{v������Åg=�x&֬>�g�W�*�L���>k*��6�:�v�O�FR�t3Ͻ�P.U|vb�����*4�l_*�lY�͋��2�i�+&\�ܵ����C����.lL�[7��5�F�dBd��mc�����}������}Z���t$���6�|E�����F$��ːQ���nF8z
X��M� �u���t�텭�����?��cr��� �wA	�S��Sl�.*.�Us5����uB�1�0<-������х@��,PA�0c	�y��X��e
�o]���q�Rˑ�_��o7�t��ɝXL7�ԋ�c~C���U����7S�/�y���G�zC2}Ė����1��F����rY��*4Vx����f�W���ɻ;���0�>CW���p;��q"�鱏�> �p�?|i���K���7�]sz�'\3�;
y_X[Y�鰿6�)ْ�����@������0V��"Pq�Iq�9�SY,��a�c��y�n���%~{�*�6%����Ju�1d��D���Q��B�\Zc	v���7Su ��J�&��b�������Ү1r��t�Bi���yMb���n�e�@�Q�	�}N��u�Pq�`Zi�v�.�����<����3K4����P'S�Y���s
�h�cA~L�]�|0���Hv�:y#��ȋ�까J�Vt�X��	zy=�Ų���=?��rǵm&�o��-��g���a��~3��� �q_u"6�}M����"ĺ�ǡ�|�1�T)����sA�DV��(�,Xʒ� 3o1�v��u��̾�o���.	3�ih�_b�X �}'�>C����8d4�9�Яzn�0/���A��'�����H�Gi{3�V�����8n�0�kY$?4b����
�n��0#�J_���h���O���Z�\ �r��i��<�Q/��[��&��-���}��
�J*�1m�E2@���/>��A-ၝ�Z���|�����i_�o��Xd��f9�]����d/��%�s���Cq%�7��R^����U<�ؙ�4R3cP���)%��}���I�!z����q{��~�뗩�⢈���\[	�~���C����@�x`�aZ���.�l-4��q���J�B���ujӘX�˦�8���(y����n��j�Κ�ʷ�<0&k5��%�yQ0�0<��B�)����������^�E�`��<�0�+�3�i���!;F&���
JQqI���7X�@������]"WS��R��O?V]�b�g h�������/�w~�.R�w/�P#�l)��>�{��َ�U�Q���l�PMd/gv��7rlؗ.����<<i��Ծ����+9��l�]�L ���>�S�g��T��/�ow� �� xoz��}��75�rq靤����J��ʀ��w>u֘���v�t3�V�`v�KSR��!�Xシ�n�*X���I����g�g	�5 �� xc�ɚ�嬥��x�*��s��V���	�����f�3�l��ᚁ �F�y)���h���n�����B~{��Sm��jť���\ e���"�v����Y���mAp�t	��;o~���W_�����׺��#&+Lm ~�6=�'6�����,_��ƯRe�;@�ʆ �v�? w�)p�ջ~�Q�M���t���<�(����)]���~�=��\v�u�9�cS�nD`M�QI��1dn�������b�`8�K�z;s��T�qR<,����u���*���XAL���{<!�;9�%�x�L������*�?�¡op��Ө�~���J]�e|�e|m���b\�$c�3�;���'����`LdE�kY�K�e����̂�O�˹��y��d����O�!e�HaH�9�	�A��~n-T6%ںhR�B|�Ǘ7��U�8�FmX�;6~���8�3���i�ha��(]`�/_�}�K�`�=�J�@ǔ�촾�6[z)�}²�~�aG�@��j�DT#��1~y��r�W3�ꏰ����R5㝗C���Z7�8&+��0�� �MF��8U8���c�F��'�Y��W�=\SK��{.n�Rfu��%Y5Me�s
#!A��!�6 ��qh+���V�gG��}������ޖ�RTS�ڏ�J	�ʋ�\�EC��y��R/���q�-U2.��LRn�&&Se�b�E��7D��-տ���X�І`%�{k?�{��O4<��Z�4���>�vC45�>ʱ��%o������ݻ'����M%#��.+n�n�E��;��w_�rB�/����7)����~n�B�ou4pF�{�t\9���.����]f+�h�����RZ�5/Vӆ�m�OW8��M�nf<��k]_̋i��4j�]�\��U����/ar[�OB��訂���뀭P���]D�m��H�^�����>5�:*�[v*�%��p���,��GyJf�iiz�:,:ʾD�"wk�|"�:���p��8��E#q�-V�q���D�&�fy��f�g�i�$)a�z�m�B��`�O�mˌ�x���e��m�J�@��t�/=�-�s�U]�:yi9~H���đF}���ub��o�LԞ��v�٘�
JO��Y�|�	�)��p�=ט�Ղu�q���+��{X�F�Q��i���� *�v�[��\�ck�J�l
:�w}��s��y+YNM/���ќ_[�mJ�2ժ�Q��ɾO^᱉�%�>R)��*�=ʫ�x��n���V��
��0�sw�7mx  -2([�N���SpqqiN��Ϫ�!�ok�.E�����y����0��eS�ϱŨ��p�:�4���7b6��(�?Y;����[zq�L.��5B|h)c�=Wgёˊ��ɆX�n+SUFaa�r�{(tI�r�0�3��ӞW�lD��q��D#V[���sX]�=+Uґ�Tu���?�uȲ�:+̈́�\ʻ���f�>�T��{��t�,�.B�J���iS��;����e�$�) H� �z�HME�
Y�.�C(m믏��=��>�_�.�
Z��>笞�!��*��ZO�pr�+Lē� q��	�FN���|\���nT�x��Sݱ"��lJ)���(�()5��+��q�hM:�r2���^G��D.�@��ʕ+����K�;_8:�R\�^){[9��/�0��y�e�:a�挧�������6��c�Șr,s,�� �ty{�\t��Da�����V	X�~R�	��C�������ue���`!!a���M.�GV����/T5E֨�t4� br%��R����,�໊R�wnp���(p�>s�Pk�$]��>=�o������*�<�0���6R��a,O�+�YU��:2S(�Yo����Ou���j���٩�*瀞ZXȫ[dڐ�K"�d�Ф���q��G�H8tG:�
�T����\|A5�BMDr�꽬���������\\���QQI���C�ȩ�=2)LRh87C9Ξ�=p��f�^��$��}Z: ^���>��F?}t���������ze�D�+�x�:��������ӧk3n��Q�~5Ō�BBB-o)��W�[i�B�����2��O]��`��T�$*iVDS���e��wsu;SQQaҐ�w��J�, :��Q8�[}����Y���?������B��]s2[3A��V�4�I�{���i<�S\�Rw�@��S��Mz�����ީ�l�8s�n���RN�.�b����̖�ȹ����}�S�}a�nCm?z3�'�b��C����!3>�K�������������nnnT44�YK@����(<���vh}8PB�SNIF�=v��(�;U-��)t%7��|�>�����T���&����q'����q_��mz�}����&�4�o��e�.ZƗv'��S��YRM��5?��C~ւ��=��P�q��-��8�%9
�#�a�����	^��Y(��8�����
ϥ8�Ja׺�t�� �!�Ps�?����'�-�#:Ԟ
�[ƷZ&�6�vW������ե{�h6LW�UI٬ekhL���9���"��mu2%99���)�.�(��q�'����� ��s���jj�j8��{=D��gHد$Q)j �v�����G�Frjj|e*nЪ�Ewv�UzB��0^����?0��C�@�^W��qwp�H(�49�`�����A�ޘf�\�H��b�֜�̱�F�z��H7+ΩꖆgK�y�Q���W;C�UL���c��"��ȉE	L��U
pf��4� ������sV(���N�揑���ǚ�r�M�#�G��YRԏ��|�W��%o߷9J̗��"���Lֶ�m�ST#���x�;�4�
����� �r�MʱݩѸ�g�SeT?���/$�wЯ���ِ0�[M�f+�*+4�DB/��C���z��ꠣ�a����d�����l/��W5�E�}wz��d�~��AJO��ً?��W��$���h�\Rf�Ђ/�m�|�k��s�E5�я���5���!K��-B���l�
��񧅖.ԧ�>,�k�Ύp�ė|��������3�I�Ӑ����|\�/Xic8�����'_������T�Ӓ[�E(m�X� �Ӽ$�(4��QͲ�����Ix��S�(�M\~����k�K�,���\���ݗ)$6�� �
�p|H)q����n��c�b�|��&;��ܻa�K��_y�/̩P�?M�ĸ��5p{��k�,�A/1*>����|��It���vh�M�_��S�{�2}�	s��'nN��95����Œ��c�|Ww>rQ��S���{y2�=��b&��W����_��r�<���8�NF>���b�>�յ�=Z�:o]�B�[�A�4J��L���՝�Czzt�D&���$R-U������������2'�~��Y�-;>W��M�������Z�O帩��+�#�Cj�y�q%�!���>��3��s��+A�=�9���\��K�@���8"��՝ e�΃��=V�up����ѳ�r񜨙㩆����ґ���V��Q~o�P����fle��4���	=}jX�*#Ø#�XRÏ�,���lFMXnou�,�Ki���[L��p��=l��j����ל�$j=P9^�R��覽13f555�+�ڛ�)���::nvW".����()u� ���
�ni���	�Ô�?>���t��]W-֐O�ޙ�p���s��e���%�F�<u-V��;�
R1�'�q�ᆯύ�ZL�t�a%�lg�h
��i�.�h��Q��џ�П(z��������%�1o���@�r���z�H?�]cz�m��GF=���$�Y���_L����XE&�#Vr��~G�ܹ�ǒ��U&�a_��[|!C˛"#O�����c�7�4 ?d렗g��QMGm
�E��#�t��7�^��V0�0���7��;avB��$(8h>�v�e�����Gx2�i>��ƞ�ta�'O�:)f��o�;��������~B`M����x���͕r&Z\�2�*_��ڌ�I��œ��9�a,��;�9��87�82�ѠW���*lҐa�+��zЛҾ��XU^L�?���Ak��n����\cv�&���zn^�li)u�r9��h�l���|nYaPZZ��<̈́����AM���#���a_=v|�+�(��k��Ž�Gx	��S��>��b�8�6��e !�D��� ����rμ|yW�.<]s����F�q��N
Vf�f�hֵ	�qVJfN<x��ėT���L^֕��Y��&��s�h��*�r{�-�殟��]7{q��1��i��XJ3�+�`�;�8w�2�|��ի�U[I_�S�tP=Ar��AK��K5���3�6�k�V/U����d凵EH�#�qϗ��ئD�X��v�A�8|���oܖ��gs��3$��ݱ�"���`�$!�{q�`������ͤeL1������y8>��"QF窝��$.A�o!�� +�:��nx�{+N˱
 &��81��O#3G_D��%��o���ߵC���$�@�ab.)�C�fc�����G�],j�Y�tw�B�����
]6��օON�[GAW�u��
8m_�ui�ŉ@�Z�����MǠ���a��|�	��_!vfSg�V�:w5̱ndLs��>��a�tyb9Y��%�%��o>���
nte��l��\,^��ؖ�豮�lPGṣ��ݠ3z�;o��|G���C�Z���y�X����<u�nX2ܝ('Yf��L��Կ���g�s%�s#����h�6F�i���E�{�Ɯ���� -o�!�v24��Q�;X*&��n�Ǽ��G��Of�I@��@1������9�M&���j$��ǻګ֌�'��Q������k�� ����TX�8,\��S(�,�Cա����o�Y�N��]�_���vUm�r�7*�_a��d,T^�G�gM U@Hsmkn���=�C�X*��AG�����"�h���сe�N��B�����Ɇ�?iCV(k����|�I�� ��X�Y����d��)�����mi��+Eӽ�=�� �=ڮ�F�����h�}6@c��r�AS)t��z#���h0�ݡN��|6�syȣ2x��gd�0LTr�)5��������K�	H�mg�J���s�,�p��Fc
�Wɲm�Ɵ)��om�"zCY��!�֋�;.;�a�.cR�X%t���e�]]�}�m��ZV�q��W|;5����9���1����J���x�;x���೙Tڟ�ԕ�Z��dG�0j��"x��A�=G4�.x�G]�Zżc��T`ӆ3ޒm|�������ug>\[mҭ�s5V���j���ԡݒ5��҈���9矷i��s�S�K� �0�NL�7f��В��B��]Ug��)6��gg���LpM=CJ��hT~�#�VG�m��X�S�!�H���
jˋ"�{�5VhM�8�l��w���j�������|��R������o���~z���[쮍s��`�C���%��Bf��P?�y���W`�5�;����c[�lf� 0b��p���Qfc�/)$�ä���B�$���fi��uS��gu��X�7׾�ϑ�x��z��E�}�����Դ�;V������C����u�"C�V*E���.ƞ4L�|�Á�[^�5#�S�m�=���l1�CɖL�.TRW~�^]R7�_��pr�g9�_.��M�K��H�>���N��R.<����hC,�c�G�4�AN� �mpii&q�'�܏%�j�	b�TTx�[M�MoDa5�f}�W*���IP����l����q��<��e���d��$�=yo�%��<D�'PX�d��&̋$���`�J��ﶔ�6���߉g3>�v�P����٨n���;��NVF"Q���ƏCʇ"����'h�藺+K!֪��s����	�{��]шJ����#7DL���ǃ��s
3&���%�|8U�<��r��Y��ܑ8��}�u0&��N��ܽ�I5{�)��[����y�4S6��[5IL��u�:h�N�.yg��NÍ��_4� t)����d��N���z�vq�d�����r<Nj��D0�h<�ӹx��Z�mF�D>�!���ق���0�6D����{���?rhFW�����4̣�e�'Gl��`��czoj�u��J���C�5ߵ�?�Ŝ��>N*�����Hy5�u�N�*u�jn���]y�ēD �����������i�)��T�[�%�� )*�g�轓SR��"i�>�4�Ј��[]�Qҵv����æ`"���B�2Yl���J��9b��%w�E��S�tJ�����=��6@Q]]}2�	��&���yA?0��3 1킌}˺�2U�X����sA%�t��)wy�֣@G�J�ab���/皨2,��u�L]62��.�M��k��{�Ez>�#��5Ţ6,��sL�cR�WQ3�]@�a)��[)L��*�z�z?zn�7�e�8)Êsk��S\l�!��f�m ��m
����Ņ�������(T��ɗ��78<��ì8��
��Au�q�8��tM�ϖ���|�Թ�>q����x���?��4�mZ���K̨�۴rz�������&��Y��O�D��4�<�'�8�Mf<H�҂�dvVt���w�pQ_���j�-h�[��s��f���]x����N+���rE������*�rc����t@ca���SLB�{B�zt��̡��ޤ	j�.\>7�,<����;��k眗 ��k��m?ǎ���&�b|p��';���՝E��Bn��*�%rZ�Z�Ň�ǐ�1����60����~m���5qZ�w��=J�x����ّ.]$�/Ƃpv��vϟ*ph|h�ܧ,�o�K��A�I��"E?� �v,�G��8��#>EDP���b���ʋp�D��9V�7<k��	SU�>4��dLAEb�Y���Q�`�����OBr GI��|)�[���Eu��R�<���f���#����ѵ�(�i�b���9�K
��sٱ3���f�۞�����lw�yl�֔xϯIVV�F����o�B�;��:ӑ�싫\C������j�Ƥ���椱��\���!໔�	*����rd��{ţ���e�'MV�v��E�s�z�� ��6)�๬�kI���PY���̜e����[#Q�^r��'�m�:�Mf%�1��G�E�� Z���;F�̂�S"ѽw˚���5����}�Bܸq�sG�
S1�m�����Eノ���@����$� C�-����$�sxX� +�}:��u�2���W>�9j�����t�u�U�օ�%y`���������5*�g�Z~`��������� �^갏W������3e��9`5�I2T, �Yv쾚 `�0��BC�����IQbb��0����h�-��|�o��Md�[6�Z��N�RXҪ>�[��D{cZM���������+���ÚC�l@J1���"Lp~<�n���%j_�e�z��쟎=(�dyl���ȼCR��� ���)�K�Q6�����>�$�{�����Ǆ^u�Z�e?��� �n_kى2	΋g9+�Db�˿�~���_��q��'���fk�>&$�O����y�s��p��6�ym_�����gvR�-���q���q��Ecm��8���Y�H�C"�a
�r)��M�X�n�'�Sn}�U�FN��+�ܛ��~���l��EX1�F��k`�i����3
O~��o=��q��	��I+�KI>v�4V���L��BK���=�[�wcE���*O�����T����bF�L�A"�dgHlI�
�h��0U\�j	�:�:�[�ob���G���S[ ��k��8�>���T����`A��=�%���_#��y"��{�ԧ�����D0߯�>ԣf;o��
y�xs�,].]�J�O�m��|R)�kl!��� ��<����3^\\��h_�Wl����]"��+��@������lоC�I_��ru��j���	�|7��`�ӛ���-V3+KRSouvu��T�4(����b�X#�r�j0�h������]]0M󷐗�F���wd(������yX�҇�D7�Lm%Àژ�D���G&| ��R��Ϋ����xx��L"�S$��0���B,�R >�z~e6m,���ur~N]�]�m����*�صԓ`_����12::+)!?a�ʁ*���AC���;}���W�[��wԆ��Wu�����U��p�xǲJB�{�[��^�~��A3?���ԋQcF�F:Uo�j����3Q3���#�h���FW0f�RU��I}�A��^i!�
-���[SHm^l���J�TW[caDn��}��8��1	4fR�yQ��1-o���*R���Y �wh�k7s�D�r6tT�O�o;S��ѹ�b�D��,wh#�m4�u�m��N<|�>�I7�O�ȡ���z/���1M��\6���s^i�ăI%!��37n��I�%v���f�4Ynk+���i��h�D��V�so�g��4+r^jI�F�DSG<��۞���?.غ���M��o�}O��k���VU�1z9��یwn`_��]W��D�ɑ-ؠQ�Dwй����F���@@��.#-�N#.��dv�А_e�	!X��Yt!ܙ���^��4!��~��#k�~T��]/@^��y� �g��Ւjr~��,����N2��n�jɾ��焚��X$�)�`n_U�x��釟cW���˽��j4:7w�ٟ�a9�%�P2B=;Ce!y�9o�>;ʿ�H�����ܑMQx�F�v
)i�u?�?f�^�_�4���e�5<�m>�a�ZHd�0�E�U,
�ؤ�-���Դ�݃Cc�5��Di�j  �j+u�J˯�ҩ�o(�G�;��U���FU(w����sa�_P��_&��sI��څ��F-�� �B�=�S�Hj���<�￹*��u�������?{�w�ֿmT���_��j�[1���<�)0�F��A����+�T������i��I�vz�g
T�3����>@�b�r5'���j��i���5E���#P����R�s����������Y�T��C!)�풇��?��gXS��7|EF, Hǂ H��q�&]����;fQ�
ҫ"M��NP��{'	���Cy�v��?Ɠ���������]�����MQ�s��Y�a��@�L�䨿��������!�n�
��E��T����� �PK�t���'p�ۅ�c��t�~ <�i����`�qd��(V��G�X��q�t���Z>�xp3M"����U	��)c�0m��qm��wWS���ܩ�N-Yoj�j���������g��?x��	���tU��چ�}����T�?4�O�W�Xw1F]��IY2L�W%_����q�7 �ם7 �8�A[�	à��s&[����6��U�>&�(����Hp��d��L�fW��e�co�n��h[k$6�~-���H)$���]S�/�����ӝq^ɑn*蛁2X|�`�d�{t��f���?�י��Vw]z8ts�i�/��7������̼����������U�?�赊%kfJ^__7��0���;)�y�Q����sf0�:a�{�]�?ə�[d͝�S2�]�݊L�9��]��˧!H��Cߠ��o�N��pY����Y~��y1#Z::�{p�?��=%M�:ːW~�*����/6�����W��@��d�����bR?�]�-�:==-���)����Z|�f?�d
v撂�=�Acw��T��q�'?}���<�@7�}�����URN��6��n$��8c��E����+��=�˹;F�a�1ێ`�^.�g��ny�:��	� y(��W��Q������ZXX���g�#��������X������WN��o���q�L<xy�C�"׵�w����P�+wZ������?���Z<����z��*ɝ�{ֱfKW[[�/�s���y�qOK#�/O6��v��e��Aq�Ax�rg��ZQ��D��bֆ�5���[�Þ�|=װ�Y�6��ɟ��_Ϭ������bv~hC=B�����g���gn+#�a�y���	9�
.�m%댻�"%�Q5^[��4ڣ�v?n�;�e:�|�>�W�,h?LW�}M���������(��r���ݻwѣ�T>აQ���5��lK��n�ܝ^ `kr���un爣�7B�������E��5ɫ�3�彛���#�T\��"�N��^��{Ù��D"U/��!��������j��LK$��'߮b�|��U8�q��6�̦��-7�L��\\\���+�em���l�z}C8�Ib��/ ����+B�����36��+s0��/�fh֌�i��+��s�8���<1��ϼ����[�g��7M�-�9�ܲ�7g�Hʨ�q7��P󱴴��v��H�R\�;[�"���L��n�1�h�6��FPc%���y�S#��\�[Ȫ�{+E��~C6�׊^�T����vÔ���cBJ4��bU���&��]a(������憂��~��%�WK�O��}��>�'�KB�<�Q5�Gx����X�O��nmp���G���D������#�C�KߴE�e1v�5��p�:���+���	���l;��Բm��ܘ+fE}<�joƻ�~�޸ULn�?�J!�7����׋Q���ޗ��᠓ɩm$��0���I�wU6�Hn��@o��t��АT
6���q�u$~���ѐ�ɞ�"}Xm�����\p�z�M؄��b��{b��pU�?��#ˉNL&�i�zs�O��J/��ܖ`�ِ�O�'��ΠZ��*]9�/2,�5�T��Ν;��}.p;�|Qxe)ǫ�	RSH�L􍫂gN�`力.�"yk�f��.����wM3��A�UDb{��t�d)�Y��7n���#T�(��N/���W�F�&�ô��jA��EF�����wWF�/�y�D�'�}}��r����O�ݻ>�q�])�����O/�c&��o߾��O;OJ� �{^�0�gj���<�HO�d�)A�ӫNw�9O� ���P����#�G�X�g9���uڸ���Aq�A�m[��_(]�ٕ%z�ș�bVF�Lʀ��MvD����J��B���%�p��1c{_is[��-7S�02˦�PA��Y�4
}H��㦡��`n�RR-ߪ�~טQ�Xyzu���S�p ��S������M4�s���	s��ѹҠ�_i���)
�0L��J�W��qmv�r��\Cz���\�˝e5�p?��T��e�ꍜ�LS=\��sI`@�6�}/4}���v�^}6
��CbY444�����BBoT��P���U��H䶰R#�	P�R��|�/ݵG�/�����V����H#�.��'Mw��-��pP���6w�}�ٶ؟]&��Z&��g�pJvw�m��-U����iҶ_	�P��j$��iMo�o���ʖ�Ni{�Q44�*��l�j?:��;�>Qc����:Cds�^��<jl��,�ZTa|�t�$���L2@QmLE�vԿ;��*�3��_\�/c	<Yy�+�}�+����C~���D�T�'N���,���bvC/��R��Fk�Y�x�^�측�Fw��b�F�K-3V���z��3`+DП�=�Q��&/��U�Mxy<Kd�q�jz�I�p��0=D�SRY?�K|o|d���?��j�J���N���b���I�п��9�F�̟8��1�����0����eb�b��d�Hg�,����� ��K?`�������`�6�� S1�'���/��x�����@���Y���㴢o�Ѣ1�V		�Q�"�h���~����z�q	g��%�&�҉}˰����$���+Rׄu<MD��!�6X���BUIA�������?�I4CڥW-�����_l�J��xO��e�ʪ��_ۍcMO�ŕ���L�#'��\Ԫ�>R^݉v�l�0~&�|Ʊ%9�ַ�Z'cj���u���n��4+���J8[i��?y��ɤ���N��n��l�c�娅;qF�{[Щ4BT����|d�S�Ў��$����l�G�ͯ��X�&2��d�R�=xY��s�	��n����%O��Hc�䇛�g*���B�Շ^ ��5ه6���N7��W}1&�N�G�tT�D�������E��_:{�C:]�ZY%V��[7G��!W��~��H���+��s��<�,�����H[A�jG���]�����y6�+=��_����Ք���^�0�5<)bSW��Uv���rcF��%�+Ȳ�����r�={�������-�9��O��E�'u���,��a�:O��b�K����%f$B
jd
�N.?�������_��ˏ��S�*B�v]�3ڳ�����k�G/%����'XX:�V�Ϗ�Z�\T[�wh��^�87c��(�3�&��+Zg\�Z�J�X�A-��@l�-m�	ſ:�߅�5��5֨�3��+
��4.�&j?�{���v:�;�0��_��J�o��*��e�Л��i�:�Ä�%���oU���y�Uصsk4��|���V00��P��*T+q)�2��n�y��D40V���ڽ
�=��*c* ���ߕ�1�eA���Z�d!M5U��r"�P&H��YE������B�{��rJ�u�����p]/�o�o��5���Vc0���5��V��HTM�k�EQ'�'��F)�gO͇�9f���],:��\������Ogъ���'Rv{���\fa[�+�����eȢSȄ�O����Xn�r�4:���%B���T�1��t��B���A7W����Ӌ����cj��C^_f���*��p����1%�@E��Ԧ-Æ���~)h���o?x���\��~��^+ n!���[ث��iUN�FI�m��M�
F�u�u�*����Һ^����#���ݥ�ZQ��=�N�f��?s���x����������>��vP�F�n����vkD��5�ӅЭ
�x��;Օ�7c���S�J���/uʠ�N̔`�*+_�(w'�4�|J��US���V&[)�Â�T��)IF����H��w�a�M�9n�t�DC�I<w&m,�eׁF�� ���	�2A��.��.]��n�j�9��
����ͩW2$��x�����؛�.�gq��o���$��V��Q
${;g*�q�3��$Y�6G���b[V��!��ԃ�� 't�7�wa�[�̶��-U{�ZV��w����l|�%�g_	re 0M�q��bW@�y�19T�P ��q��%/riL�Nڊо9�qg���[M�]�3���"	��W�c�m4[v;�@PK��-F>Pz3j�4� 1�����"Y"�t @�� mTG�7H� ��s3eisI�}zQ���^�
ڐӳ��a�3�qa�b��V�����75_�m֟�ON�/��n�u��^��V�h�R�v�&���$��tf������R�X�	M�00�?!͹'����!��#>����p�>��p+�LO�ן�ɮ"�,^9���k�ra���3����ֵ�nkC^���3ˬ��)� *~�i�
IݮN�p���¤�I>��(���B�j��,�E�M4X5P���Kش�E���ӷ�:�;�8U�)��)mw��s��_}��:�n5K�A�{��,�$��z�A�?�6uƐ��hY:B*�;�_�O�n�m�� ���Y���WՀ^���;�U�.��Q�o�L-8\	KHtʸ��t���d�B¯s ��̪��	��Ze tƩ�$���Z c��yHRdɐ���/cǊ����+Ɂj����.�G�}	�����}��ص	Ξ3�ޟ8�ݦNVV�d�B��̊�K��笗m<� vNi$CJ�ތ`�"��A�L�z�n�L6���_��-��yb�b[��@R!�D!�������N�iI�qY�o^�]MM�&��1B�ܕ	S����K��`�D@Q.��I�"�9n�5��VJn/�Jb+$L^�n=GO�(���eT�s���S��or;������jv�z?	�?e����� B>�艍�MXƠU�G�k\�ՊV��Bڮ�b�P`i��SK�y��v����~�;��Ʋ����~�\�m]�97#`��c�%��}�u��	u�F����f�[wZ/��W#9�W����xz���r�S.r&	rrrBje#@+N�Y��%�?� ����K���0L~z�V�!'�T�"��toXR�8/�9��Oa����H'S��_V;@6��T۬�V�Q7���t�"�:fp.u���._茇o�Ɣ�����n�,	�B�#��E�U׃�
߸�l�񽒜��3﹯��
���.q6���KW|u4~�_Q�?$����]`����:�Pς��;����a��B|�X��,��O��s"ތ���?%In洇?����OpE^v���1�+n��	1G��l^�6@����g�υ���et�Cvr�*bТ�S�j,�!�s�j&kޑ���3�k ��L��ZU����H�u�.5�I�1�P� ��e��h�������ϡ-T<��7���s.X����~,�Dw�d)�|���6}�כ�$���uk��Ҟ���X�ʲ�$h�Hx	�҉ JC�ъjjnʜ�IXt�Ĉz��a ���>3���{=[���)�h�Zۃ��I���
���
�ޫ���s+�nA����J�lja�r1^{��o�˗`[�q��E=�1k�{F�ZHO���Q��s���Ak��U���sM��{j &��,��ĭ��(a]� གྷ�Z���}��OY����S�8NԬ�����R��T/����k�
T�ɒ�W�j+|��k�v������W[�z��z|Ǟ�R���;�ށG���Sf�' 	���ِ�ʇ��<&$wXD�d�v�*�z��id�R;�����y���-�G]�Ɏ��t%[��&���6�K s��j�v�է�GgńQvU3��3��e/M��/D��yFw����۔�c�M�n3�Vg�٣��S�2����'��Z�/0��.�IO��р�$;�_[������հ��]����F*6=�&��E;rU-1�F�[�W�A[��j�~ޠw-4�q�� �gWW��N�aT���Ql�6L����H^Y���ȹ�V��`�S������W�(���yR)XVdX�R���}3/�G�((Ft�s�;�ա��{�e�E&-T�Ɯΰ�zf3��U���;������U�5���?,����܍-�v��G���y�|�q���w�4=�"��
; ] ��d��ОS<;��wWG����K�Ә-?�����e��D�#O�f�3��CT���@�$LvW���:d�N&���������>c�>~A��74�'�`�N���{��|)�9D��gn�D�v�I����a����HX���5���h�DT�F��A*���p���� �8�8��_����P5(����U���K��G��o��[�>x��8J���flc�/�2�Jne�8�r�^�5e��*_��Du�g'�s��ŏ"[���\o/w?S�T �-~XQ@B�������!au`�ps*�Q�D����X�,���8�w�g_"�3I,��>&��4҈;�C��1_���*�B�ؘ2;���)-��=�HD@�6G���cB|��.=��?��B�8����>h�b�
�|�3�>���7fcjm�z�/4���㗤s+�ݲ���dBm���s�=;~��W埠�y����m͖T�<L�_N��7+��vЎ|�:���]+�E/t,k�a����>"w��|jL��I,�r k�?��$�0n���-"��`��4Qz�w"W��\zs�&��c�KHH�&]�&Y�/���HZ�	:w�Ŕx�V̇x8c�1�zN[����#F+��zE�5<�o� �i�m���m^?u&��8a�%��FQ-�)����NrC �M�B����Zu枥�v��_�!�P�(�a�7k�7nf����d����^)	���
3��*�W�Q����a����
"�q$A�.��~�WU��td�z�'�l� �y�U|�a�>�����Mp媧�C]�Vb\)��Υ�����P��`t8׋��=a��8���F�x1�������o�LZd'�é#i���қTYۛoľ���%yԉjI�Z(�����`M)oV0[e j�o�Gjq��<L~�/TC�N ��Ԗ0�ݴH��r�7�l�D}e�k�1l��K� %���!f6N���k~�i��9�����ˀ��� ��I:F�
�6�ƺ�9�lX���P����~3��YE�3m�]A�^���`Vv��W+z����'�������ͭ����N��v���}W��>�O����G.�P�ao�p�{_��^o��@���D{Ƥ�ki�Qe���惪6�]$���ЏU'ǭ�)Ab�:�Z�����|�zt�����S�����2�uCVd��<5>�SjF���^�K�����D.�Mi"�&rB��4PuN��K��W�q�` ���H񒻐��X�?x���-Z��Xc^M�u�@j�A�W;CCe�2��g�7H�9���gW�_P�B����]�44��'o��~V��8���9�e����}�0�B�㠗�+|כ�13Gj�Y�$W�}�p���Д�Y{����^�
�j	���v�eBg�_����Y$}3�ؿ�઼]Z���C�S�#��n��͆�s���a��l�Ķ����� 7�.θ�j�%�"@njP�	fr�ns:"�%zC�s�����jIZ����^�֘����'��m�z���S��2�q��%���2���F��'gZ��S��A嘏�wc� ��v#>����A�.̖�S�Qn�t�Q#��<�����t:�N�VhV
��mX���j=˫b�a�}����p�M��|�L9���s����%kf�F�{�*�����V6�t��1;���p�H��X|C����l��I�%���u�r����:��Sh�|�Jn_���{�}��eB7fL`"$bGZLj,�J���yrw�o��e�W�K,��r�~ۮ�0{��g������VMdd�Űz}��f�
%f#�y���ȅ�LճIǎ/z>��Cc[}b����)�U8�����6���F@S�[.\�OƂ��&����Gb5tM��v�ʲb��۬���Z�i�)e���ug�ACBx�	P�?���OMu|V[p��;ɨ��դ{)�&�1�6N`c0�Nj[��[���5�>��]�X�X��l�Ns�+����;�����U�I�*�O�����;"��;�AyѮ��7��V���b�G�A�� �F]\���}��J�s��`}��H?&���2Ȏ.��]�t�َluEd� ��k�t#5#�g%�� �����:�:1��
0E~t͝�N�L���`è8!�j�� �2�"�v��O�Mp>�vI���`���)��#����5��00�kw�{ht$�?�\��Z?O<�9����c�=��Z��9ʑ�홴�m�%�j1l����L�15�´(�[�CwK/���J��Y�UKZ����F���;�2�L;�֋n� ުA��I�3�Iw�������tu�e]��B�w�g�
9�:�H��lѼ��U��ɧ���ϩ��y��럪?��OZ�{�R\�Oq�t�꽠��n&}}6@�e��Nj(��v��B>��LRK� K�[��5�_�^��.�I�E��#j$���W���l����O��)���WɆ�l��
S�����>��_�{+#X�X`��p��,�u�u��)ޕ-�؉���Jg���o���r^�k��e�ο�Vyby�]�j� kQ6�}�[��9���d����ԊcĆ]��}w^1?{7�}����,c6��`'�P�Q4#أVu26vl S�-*$^�S��'`���c�m燧��y��Ђ����������G,���=Y8V��?Փ��/1ozQ��l�5�G�^L��&~-ɤ��#>��V���n$}Ό��=�৿�T.�g6 �c`)��b�(qxXg�1+E�K��6�E0pTB�W.Y���7A3�{�L��aa�
��9躵0�S>i8�M";V�#�t��CK�շ=��f�ӟuP�S�r�=����7A�������s�fP�)�<��M�x��7@�ط��eF�s�g��@	L;�4�Za�N4\�<F�(�+���W&�voMd0��hX�H�F�lٖ?h$Ȉ��j_��#�������L���Ͼ��ghⷁA�O�,�)p��e�lv��e�M�IT������Q�8I��6niG�h���j�`E�ט��B�B�� �?�3e��{�k�����ì����|��F{�I��a�`_q���U_�;��Џ���������K�xg�^��! V�U²�T�F��*�"WY۹6��#)��32�l���=-#���no��j���W�g8X}L�h�n.�؟�!p������Y>��W?;ҞX����W��r]�~�K-��'������U� ݀�����c��*�Q���������DMy͸J8���2�\�,���=��ZS�� �?����B0'�5����r�+�X�Yd1�ܼ�w�V�[�j��=Y.m	ׅj���C�@u4�wbL�%��OL%�NA�UJ+���� Rz�1yx�������/f�2��,{?��lw�\b2qt�K{Aa�u}�c)$��U��P�iI4�6F9�������H���sKz�ʶ&��5�TB�VR>rdG	���f��w��SVy�-�U/��\}��_��Zl7V(�P�i_�0��J�����k^#{�S��e�@�yGۿ���L�-�̄ĶT���a�HP�ip����hZ�EO��	"N�S��ٞ���Rwr��g���ʹ�͚���%�5V,i�ԙw^�2/p:��/;paǻ�Q�������m���ۅ��+ hp]��,��ov�� h���or��(�0��ON���}��^�3A#�w�}�ޏ���u �|S�d���%��=���R��(���|�V��y�qN�,����ν�Zz4<�ϣ���r��b�����Ƭ��{V�� @<R�	ҫC�F����Z?�7�0O�״d�^?���Vc?fE
�"W9�X�奕=P����C[6j�I�*�$o��}F ���=(�Xۿ�a2�^+U�^s+�7P��S��w�;����W�0L��V��Bu�x�|�b���c2�\&�^�w���}^�,u/4��3�;K~��M=�$̱���U>pS�+v{6XAl�4�� ������0���:nM�@�X�5Z���ȹ��=O���n��[\ZB��5���3�ɺ�W����7�n8�BQ���AGbd�������SC4�9�3~��[N�tX]]��e��H�� �&�YY����$8=�fZ��_6��l�Ĝ��C����;-n7�yJ�N���sy��p�\8�N���G�G���Q�2��]�Iu>���}�١X�p��c�ܠ�����L��R����R�7�߼%���M���'�C_��9��'f���XL�~#Ʃ��������J�G���戀�N�q:�V�;w�j<N*G������[q�Nj�s��?�[���)�yg�@���@��S�9��^�VC�E�K�Pv
��6?�Z��Z��+c�<DU-w��?���S`�MdJO��8kj��5���℃='V�A�[�������!19��W|�[:X�P\��+����4�C���#(�k�l�[܂��vD����4�#�R9#��&F�fR��%�kj����r�����"��E�B�gꔀy�넬�w��k��� #C��c1����*,�M�(�զ53@F���nϗ).����+����{��`��ӡdc%|ަRz��9�/�XoO$�vhn�����J1�ޏ��p8�ӿ��W��R&FK�l�W�zt��$A�4�"���?�Z��Pa�\?�-y!u�U�o#C�KH�л䁔%�]߈ў|������J��E��p��Qn�)4s�]�u�0 �5����p3�|�:tA�Y= �S�3]���qo����<Ԅ�/��H�׎�߃W���^�7�Om�w�{����?�-�o��r����ف���;�aZ���	�@������5.Ǩ��w��#�u��;��K�/�Y��t��ne�Dv��"�:�$GX��MI�>F���ɰ���HU�B+���ݸt*����]�6�%o�HvrUB|6YB��f��ú]Y��r~ނဘEp�+=	eдO�����1�4�c���T��r�ҀYp�C8�!J�%.�l�U���cy�3��F�>jih�!�c�o�����@�?-��O\\�;X��η-r;�;�l�a\2���}�fA/J��bU�苏�G�M�3b~�F��f���ǹ;s�J��M�.��w��8Cd��ʈ���)3�&���C~���h+��9M� <��2D��ӣ���j�S��(�9a]�L9jXjj�V-3����ډ������_�յ	u@&	8��bM��zߐ}�Z����gb9 ���>l�yr�e�KjR��+y��m�>
7�����?�َ�:a�� �ESG�� ڭ�lL
A�Fk�$_�h�x�B1���j2ѿ��4��`:��9����0(<Lo��[�	�}��k��AY摽�3�E���6Lyͨ�z�+0�E���� �\�a�U�ѫa4s���khՕE�'T�8��s�]��������!�)s޲7�o�]���z�Si�"���
u�y��	�$�-m���� (�� Ex�� ���:�P����tD0%O.x��)��!_�Wd�z^诣[z��'ٻ�ȓ�	v�J�����kO(3�B�w6����vC�o�m%!S�.���|T��[�A�E�L5Xk[�#Ϸ��fb0��ˇ�r�m�r�PN^P�%��xr���ʎCP�_���<�u��v��+d����������	�+�S���l�l��ׯ�UY�3o�B��:��,6똠���J�X�i���;��u�:g!9t|	� NɊ���{�C�t4�
��̕��/K���o�W4�vQ���Z���n��������`�YG�Ot�I���xH��eOn��0f�2Q�!���OD��P4���ǥ�����3~H2���ú�|jL5����.����8���Q�Eo��@�D�x4�������<�]Ԑs��3��`�c��w����;��v����,��'s�c
�h��~2�O�ؠ�S��#�F��mFF�S�R��?y��B>$���NNjP���ÌƖ��T�jR���q��Y-Ojg�&_J~X�wɫ�]:�V��������h�'�y�I�����ִ����'�o�Q[C\�A��whϋ=2j��6qro���q�pK��_�̙ň��J��wgR���D�4	�Ӯa��a7*{�`qm�K�)K�����~�!6���q"���i�k���*�Z�e�*3oo��;�K�t*��?q�>&�;_}6�6���vEd�9���u�[�״��6#��;�.~(�Ѷ���-���R�o!�mc�dp5�=�@/�˛�� ��p^<����2�]Ж�V��+�*��?�ǀ�??��K���N�?�IT8U��=_j����5�	:�l�������U�3J��pU�)O���0�..D��z_�O����vQ�bR�A4�:5�v������^���:;~��޿c�S���ҫ;i#�?�%zk�,9uK��h"�ny��m�Ь��i2Tz�"�Z��x~��s+�;@� �t��Ν�u�.���;���;���d�v-sD�K5�Չ'=�L�d���\�3t����L,���ѳ��P�{�Y4M'{��09�<~XiZ�}t �̭�-�����ju�@��v��������6a��Q�����)h��b��3fˏ��2�58nq��A�NA�������*�̺o������PS�PԎ�,j��������f��;4�T��nT������+U`�HT���Ci=
��mc���=����g�����"���6���»���>�8�l�q��a��� ��*�7��)��*edy�$�o��|Vl���kuEh喣�����i���>�d7����ѵ����fC�j�u�GR�VL��U��-����)@$���J��l�F�lf�Ȯ�\\p��ZO\��h ��x��	C�$��*�!^�o�
��nʋ�U�tΖ�!c���]AKK�mL�[��ڵa�<lQ��)�}��Rc�|#T��k{~xjk���s��i���~��Xưh�31ә�9��N��ku�#a������aiYi��Hc���ǗF$�#��#�m5E�mh7:�����FY)B���a&�KY:�7���?l[���&�Fث/��+6˕/Y#�W���7Q0<3!�tuGQd��%T%`)=[v�]4(,�Y�y�Zr��9��c���'���������5aS_i�A��egFj�=�a��y����Kk�;>W����Y�-r���d�T}�u,tT�o�v\�qfut��yw����Q|������}ǉ>� %�|�\ {�2w�
)�C�)�L��,3�"$L`�Pe��	U���������('y��.��tdm�al |�K�ɋ����<U��j������9{��3��� c�����P'T��9��Z���u:U>}N�p��K���#���u�'�>aF_b�2(��\3*�N��5��z����,�*@+�?��C�X17ew���l����5��8���y'�(?�E�O���{�t��:���O�Bq�__����%u�׽�E ��^��0C����k��6��})���W�E+̜�f�7�2�C���ǘ��&Ked�u�So�&��%��j3m�JJ>��a�ms���W��L
��8jR�N�����>���7��u�S\��m��� �.�d6�oB����&W�>�s?CL$d�.�EƇ�)�~�!G! ��ݵ��͘%E��f��]7�z
�{%����=e95}��R��u�H��Z�s6,u�7*�|�<�"
lP�3s�C����#�1�^�`�a�4��=.½�eՎ	:�c����i3�n�&��ۄ�x�1Z%]
�ž4$%tȖ9ER���,?��T��ѳ:}�6�s����R#l,����vj��tZ�D�k�e�a�}�T���!hc��0��J��	^���/j����4��FjH����3K�i�*�mH��ҚcCwj��:�3r�˜!Q��M��>���v��fb�v�-o�l��Y2�\�,�<W��e�Ѭ6[s��V˩�11�4t�$��K���EL&P�*V*�?e�F����Gq;}L G'�mE\ʗ�u0�v�_��zA�ݒ~<�X�(>�x��w,�������Z�p�N���_�C�8L˚ES%A�w�j6�f���1�	{p���r4H�;��En����|��<�R�����*�����a4�ǅ����ɃV92I�p�=1L.��k�� ����'��P,*Z��m�Lt������-�A7�'��-ƒٶ6b�����<�����ٯR��x/�w*@re�7��3-�m���]%#_o�9q�k�C���j�3ý��Ɔc�)�Ŷ�G�O�ξ�����y�,i�{���}�u�/x"߁����F${�h/L���������?/�(�P�� 3�ۻuR�ոG���v�˪y��o�`���h���Kq��[�D+�;j^��4;r���D�@;N'Ge)(H�ˁb�0��y�B���r� ���t���m�O��*��?ܶ{E��a4U���V�Z�FI��z�U���m��rw�(|ܷX�rl�e�c���v��vZ1le���u�B��)�F���2�$*�d�L��Tc��YҊo�f���SW����A�Rh����++������(t���A��5�j	o�ba��-'6�Đ"��S����s�����U�-%��W �D�>�fG�`��]�BN�eC{���v�=g�B�^���B� �S�Σ+�/�J�s�|)���cD�	C�����9���a�G��]������O���U�A��ɏ�{+gMc1��U9��|�����߯�~4=$q��=���ȋa���<Qٝg�5��U��a�;�B~�7#b�Ҍ���tМ��
�T�Ӡ��h�LYPa�x@*o�D�5_������M�����j)�:up�L�o�x�=1ʑ5��zS�A>�^t���;K	�a7��C������K�y��sm0��K� {�9 )�{��������Sbt��~�j�v��54��������Yȡ�n�pw|l�U��{���2h���lw�o�&+��g��z�d@@����Q���㦩E^;�G<����q�ӿϓ~``���پ�F���ڗ6�W+U�
;wVΏ��P-�}1S�XU?�#��2<Q���
O���-�/얺ڣ�+��m�5�BF-���[C���E��U�US[#��W;�h��	��y��m�
�,���ڕWH�Kx~�}X���eE�K���/��JeFP��~ZZn/���;Ƿ�@vUY�/U�,T��d.ՠ6�0�~C��P��ѿ��`�"�L~��Mt��if)877W�v�������	s������GԂ��pfE���À9���c�ӟ��W)��\��j�(���{:�x�
�skƖ%�5�R��p��n��q��F��\/��o�3��I�+6�n/>��� UB+�׶�l"�{�w%�>�3���:jj3+����
��Y0�u���Q=)Y��ɔ��|�v��K���ӥ+ݬ���I棫�g/���������x��˯[#�#���F�'&<��K�yo��߄�{Q;�1� ���D2�H�v����l��Wo������[c@�w�o:�_���dr+a8�{D���5�j�����'6��� ���ax,�k%�6cX���9919�A;A�7���'��:���59�ɽ)��a�3gvl�Psu�=X���HvbY�e݁L���_��/v�Ƹ���>��m?��)���{��t�c�
���?��Ark�__�S���1��V�>io�E۷w��H��T<�v�/o��`�G ��t �M;��kp2C�Ҕ�`'q�hɞV��B�,��Y>�l���bHX����f�����t����S�m�ʒ�z�S�����4��_��g�ߺ�������~�(̅s����%�g/� �D�N߅�{����mY�N�t��� ʡ$y�������v�����@�эl�{�6��xW�ijmm�]厐�ŋ�����ɏO S�/xM��@�̮������A`kkɰ���$��9��HK�C���f8fl�r�<�͆jy�=X�l;�y��w6Z�a���f-���9�j]�_�t��ܗ�K�['���̨��Lq�|e�R�I|X7���B���T?:��"܅�î��S8��~���w��%�u����YК\Y��m-\��	(<ˢ�_J�>��n��Cy�*��0ӡ�X~�V+= �G"����ɿ�����@x�0e�I�������i����q�k^�%S��z~�=�j� �}�%���t������_l��p�sr�P.����;4�0WȒ �_�r��[?Rc���V��Wdx�=]�J�8���9��b�<Ֆ�|���s�2�pߋ|���r�nޯ�l߉�+q-��&��G�X���B|���>0�fZV�ٌR��ӿ��ph0��F�����&�$C����1��L;k�alr^ME�Wq�H�f {a��Ҕ?��WA��Cҝe�Nܹ�x�ge�o�7��~>�����g��6����k,2�]�"e�{�{!=�#̝��q?B� �*܍��L)��`^��"I���Dԟ�����]߾��Ҭmn�
��E��Er;^�Y|�N���+�x�V�<&������ں�
���ν�R&&&Ie�	�o~}�`n�;������N�s:�x��.���b�\},E���얥�����?<1#{����?�h���:�L��K�N����_GG*�����M!���R%d��Y�ڃW���؄e�$f�����;'��bF�^�W�V���$��ꯇ�[���:e�:4��hm����L��[���}C�l.cZ!���5��[F5�e�Z����\��'��nמJ  �x��R��VRE�ČcG�׺]^���y:2�h�`C����>n*LB�j�N^�e;P�Žg��gM�A�xP�I���Vcn��/߽i:�.�P.��`�.0��3{�5ɋ�ݫ077q�c��{/�T7�����:C��xS��J^��J��Ҽ�/�pN��u���[[�4�Т̫;i����D\�4vj�.�5��qF����~X�������ގ:��fh����3�B��x�?�;]8{W.�������<����ޑ�F>%�h̓F�U\RO����;7/-����jB���sF;C�P�~4�2�����ϐ`��	4B�ܸ�&�����4�N(_���`��yo�P�^D�CQ���6��"���=��rT�c\��k��Q?K�{@S�F_�Cg?L?�Lu��'h#���z�����P9�- ��]�ޗ�$g�{l���Z�����6�(N�3�9 );wIjW? p*Y�{�*J��|iQ���<���У�U����i2�%d0����0���?�����;��	?��79|{�cb����\� �����G�#�c�E�u��:�g���V�b#�KȪy�r�E7x���nW$[ ��i�O��������R�C�_�T��g��ɺ�~�v�� M�[��g^��3�dJ́���@?ϡ%6@c���@����rr�ޘZ��;�?;F�����҇Ǐ��ϝ�|��?����l�d�5f �����..)qb����(��[b�$��͖� 'i���E��p���񙇞��t
���0�������R����k_���}�����JwwzI	i�.G@@�1 �A�C��nP�kh��wo)(|���^k��x���&���݃���hw�W��j����"=�%M�"�|v��M4)Z�k�	oc��?~$����ct������a�D--XH$gDR�$3�Y��w���ޗg$�b�}�g<�R�-
ߘ�������:^�Uh�������2Rߧ�|扦���	ڰ́��{_rd���'��bœq_�8:�.C"��~F�����r��QP�0��f!�Ԙ����h���=[t���[���=@�������b������@��\A�Sg��P�6��I�
8
�	2"�:R������
�^���M�R��~n�ۛ�(ݕhF읿>�qC�k����blZ�3�?$^�"�V�X�l�kH��A�l=��&�6[4=c�_�ܧA�jy-o��X&�]��9�5��('#R�NΧ���1�
�;�q�;eX5�&߬s����B�����u��T�L�ݠ0Æ��^�⮶�}&c���|�;r���wx���xd?��P�J�1�]��:������Jb���U_1q�D|��q~`��c��=�"��kK���7�������8�}�*[T�e:�3Ͼև��+ }��Q;*���w�e�F�Q��x.P�㔢��ã�����®�P���6X��	}�"������-K������
�����K$�WoA�U��_n0{+㡳�����z�ڽ�"�A%[3"�W$I½��N���JJ=�/M�Xs�Բ�ڍd߀;�y%�,�&�2���	�%GV������+v�dڠ�̲ʧz�����A�9��:�Ѐ���$z|es�)��ƹ�����K�z�<�6�I\�qH�������*:dk��t��M�"SF�_+v}�E���L;C��R���
'���9+��qϡ��HIƶ}<��/^�bt�445��p:NR��`3��P�������h0��DAS�%�ѱ�W�_*���RK(s��f��������I�Z��f�ծ�����58�I/�����e
a?dr+	�(���X�c����u��L�\�,���ϖ6�2?]d�A���C��垹:"�$�}o���`��J��B_�X4�z�r%�F�7�}�_=�!>xtR�w�S�R,6���!;e�Ca�K��^����P��볅�`��?�z�⢰:?,�Y�);��:�eE�V���X��8m�
H�f�J�i�e�M��ÅD������6���K/�j������+cdX��]���ӝ��R&+�*�h�K���j��(���om2�)�r�{�}���'�wj*X=:-��������0s�r����i�Y8')�X��W�@�cp��U:V(�0����ՙvF���T1i��%I����̂�F�U��	5S�d C_�w��t;xI�e�v��y������]5��.�7�t-�:�"�)C���H���wX�W@Đ���7 9�VqI���QE���8.�=���9��ۀ�{���*&��T����/(=4��g,� 5Y
��V����NY���<ǃ��� "Bٮ�`�]余�)�?N��O�|���cl�Z����`�nZ�Nv���$���-�5�qOYJ(���`-����>W 0������ܓ���>@ͣ���Gzm2(j�
�,��R�e�%�J&�?�q�c�}���@-��h��p�[Vl��.qg��hΑ-���6�S'�������B�w�z �3�6c�0wr����Lkg�7�Ռ��!�nٔ���Edm\@��!���5�L(ڏH�����c��A�C�%Pp�(D�+�Dh�H��#�y��zb�ٙ�+��D����B��w0��Y}f�Ԣ���pˑZr�=R�P r�Ғ񂓑�<'OK�lD2̮U���к/�DY�DaU9����O�u�t���� �v�����;Ipp�[�I!����ZH�N�f��b��@�������5���>����+�aI�窫P+��M�X� ���Ǖ]BB�]Y���iՍ�&�b�f��᥾^�����Ó����|�bw��썇"B�r`���(�4M��&OdOE��Я�D��@p!`����:bP�Uf�xc�?q��rMII15���r�;�J���4���Q�)'	.]���7�D�d�wZ	2���=ꭷ�'��K3^e�Q}r��e��;��E���M����+#�<̭����n�R�r�ƈ��$~ZY��h�~�q]{��d��О��{��{aߩ�>��G�lv�]��U�iv)�����{�m���=)����$	 vvvT�*du�\٩����+n� 6�@�"��2j썅����Lσ֙��`4�W�x!S}��+�6C<��,>�v"%�30%�����-=(E�T� {�8nV���e���tG92@����
��ʈ�_�M�`Yڛ���J�"{zx���^���w�{�@ʿa<��Kj��� ;�k�ϼC8�R��,�:bd��^�>���Y��&F��C�z���N�Wb2��e���.���q����N'�\0p.@���E%|����E4(L	��E��<����h�ȴ���̔ߘ�t(�!Y�F6�%S=E��G��<�D3�8�@���k�T�G9���f�m���Z�&~Gq����@!0�{DjV}9����D5���>�8|>[{��p����o	@b����(/5���etר`j����y�̀
'�cT)~�y�6�����\����U]��CƝJJJ���$ѹ���ȯL�<��tX|�]��-੕�v�ߎfe1id]�V�=����Q�*�S�����|@}8���G����R���hh<����G�x��+�F�Ӷ%h�]7���ςk�[�?�K�����f@�����	��i�,#�(=�`�n���/��,��>s8�%|�-fP��!�z�H&���4�4��ܷT? ������G�B��oqZ=�'�:�k�OrQ�SE�n�x3z��!�r&�5���Aa�xM���s�/	L`�M�J�+/,U7�b�� Ѐ@L;}��mΣ��!��Yڝ��
mh��
����!e�^��0��HMM}_PP��� ͩ�1b744|w?�HQV$Jdiusp���ә��2�n`�X{@�6�7���Tт'n;~����c�� �c���ci~�o�d�7��D��tMi�l��|Se�7��]���͹��{�RK�(����L^�n��-ZZZ�**�6�oH��2H��nM�48^z�7����xL'��0E��GI��蓘����HJ���M��\~��{�� �d:،f����)�S~��M�կ�Y�nX⟄)�W�nrss{��jy��Uz�n�E���(6z_V$���{�9r���� �wn~$�)����>�=R�=���-�q���~5�S�A#����^���~���8 �vG�NN\���+�^y���e)$��p�`�����=ky�o����zz��W-(�1kCҲ߲�,�V%5p!φ�%���mE���я)پ	(��xt4ߠ��l�t@A�����BOjyO���Ȗ�`��m!��{��!"_@��R�~]�=�yߢ�?*�HƘ2������5���
�ˉ������Ὧ����P��u���I�&�M+}/V��(}(�@wV���݀e����z̏�TleO����iH�[�2���i�b<Kh�vm�C �S�=�,��ˀ�х���D�E��_S��:� �X�CHytYJKr���d��P�S1Eyu�;��Ç��W�m��64{�ۘ-P���*[ZZ���ƛ�`o{�R����«E�#��3+}k�W���,�Tm�}]H�8�Iż�{���92/����7莽opP��Lr�~���!�[���פ(3�ST�a))o��N���5WW��`��z:ӂ	��Vh	�.�@xWŲ�4����/?"�Xhom	�����R��*�KL�-�6�E/�%}�O�Ԇ�*hj�T��@���g�2kRU�J�_z\OC��.$RRB��]v����#���H>c��)mn��9�)�o�TJ��z�-�B��c�֋��a{mٟ �=U�t��o���Q302�}	ֱ2�{g@�M��^"���p�Q�a��:�}�ԇY�ލ.�1�a�A��<6(Fx����Z'�\��"�g�����u|ևi��J��/~G�9�Z���J�f�qӚ��?^��.���t�?�S����a�~_0�f��P\A	@}���Fr�Z��ֽ��vWZ�M�P4�Z6�16�b��)��Tj�(I�g��<s.����%m9�^*�V@�ϑ��C(R��Zi���.�����Tg��ER� V��_n㯭�9�&�	jT"%�=�_>�z;��	�@��"h��0�����Y����C):��P����3����F~qp�T����?�T��U�����茚ø�W��P���L-��W���y��r���fn�ڣMͱ�:��Kk9��0m����ʯg��l�����+D��[�鵻�ĭ��7 ���ߡ��e�'�P��|�r�]i��D�������o"v��Tg�yv S�~.u�s���Њ�H@����
Q��Prb]S�n�����Wy��ȵ���?����d�J�z�+E0,�����Ç��O'���̇g85TjOeM6�g�T�n}[����E�R�k���c$���ec�G�+
ëd��|���*tԲH]AX~�=!��}+'وPʱE{1�؏�/���ϣ��e�Ԋ�h�I�
�l�U5E�s_�<"h� ;hnMe辇�E;��ѭT�5I��ϴЭG�ٙ~��>x}�	�#t}�өŭ�*4���k�Xw.��;>���
/�p��_*�n�7��]�Q��N~����|(���PA(&Q����w|1�n���㨏���gz�Rq��
�
��l4�:Û�7�eF��E�ɐ���7�;���G�}����TѠ��e����x	���p���#K��	��r&���-|C$i����<�t��O n" "��1����@1�����
�c>올}���Ľ���:	ɝC��I�5���@GET6wҺ��9r�XǮmJ�꣌��˗�{�f�Ƶxo��#�����*�������Yk���R�����U5q��R�
/�Ө%##�`����`�z\���݂EKZ�O6D�lu!L�M��V$����x�CT֠�����6V6��������$���s��у�	�������a�k�O��r�ѴyBo4X���>���!���7���[H���m��~����k�ߓF�-
R� ���ǶAE��T��?9�ؐ[�z�w����̘]<<������X���_?���T�.���-nn :��i&H��&�xkS�"dq=����B�^0�5�	iP����1�o��>�����k�]]��ͅ�m�{X�Z�+'<�R��GZN
����ށA��om����OL�*{�;&؃�ԙ�������Ap����rA"s"9c:a<{Q�}_�쬕�0�~ҫ�0�(�8F��~q����� #�I�!�����e꥜>V��~8�b/	of)�á\�|�~��䉾}<�>�Ӭ�� ��v���ɁK����J8��O�NMͻk G��#��tG����#KO`��
��Q���by��p��Ԓ���uE��a?=Ռ�b�{O%~�[Zǟ��
�`_6_��#�̣4�HuB�v��:�-�����+|��+�~��������o��/7=���:<P���)��Ii��Pǭ������6��?lD�w��w�A�Wrk'. �NLa��Dm����թ�K|�}���2�F���4p�mK[b������K�:M��(� :���"9����F��7�Y���7��)�����Z��7�ޔ$?�#�����f�����e)��2�3��Z�y�Q��1����ޅ�����[���?���u�p�5-S 3#}'_�M���8?���waa�ws�V�KMv����b23[[�蒌nh]�x��,�O��;�RN2�-�N7'�VB
�
6w[E����5��/'�nb�c����4c����Z�V�j��~�6hƤ6!��N˿b� �&�[0���PNQ\{!��c���6�v�ފ���5Ķ����3��x�AAAAgxRy\%Jō��v�������Z�SVG"�
7,��"��E��C��Uￓ`�� ��7ʾ�l;P#J溽�r��_;��o���]�W76��˨��;���}J�Ԏ�J�Ԏ2X�(:���Sό"��'���& �/L �l�=t��6rsε�$Eh��Uƺ?{�����7�Ox�Lf��g��F5�ǣ��l2�Q������| � (��)���Oc�џp����p��R!��|����9�U��ڵɚ)��i��/Sx�s�R�g�M>��\h�Kw`��8�i4�˹U�A�u����sҊƻя�Ǘ��A�����K���s�7$�=Gw�Z�8��W�Ο��+]�k�$#"���x�	��3kδ
�-\�5A�ta�3o�v���`�������9���Qy�cN�tx��n��>�	@���N�
v1�l_"D�B���x�|4��V>n�Ί!E�y�Ԝ���kLfM��/���K��C�ԧ�f�:f���"I�5���!��B��x�Nþ3Ê{A&r��C���:W�[kICEy ���S)Gw�Wܨ�����#�U�I�7���G�9F،�G��T;���4��}���좛�8��&��Azd��H5L���TNR����g��������E�XQ��V�I}��B����:�r�%�Y��A����ӷ��*�x|�K�l#N#W��1��t}E�¦-b�в�k��O��;�Z�����!^�`�?]Tm�$�DP�z5xS���RX�ey_����˅�-屪�,��4�(�Q��_��ZBl!(�9͎���;�OLq�K� �~�� ��S��mP�<4l��h��Ol���O�A���Y+�x����/��(���^i�.�> %��և��4���L�	�EtRA����X<\mX�I0I�(��7��o�+g�
��|oS��җ͏���H0/�Ν
G�b?�8�����HA��O1�g������x�y��'W��"ܵ�Xh�U�UQ)�2JMo��(3�ww#vv�cx�f	��Z��,�,-��Lf�	���RYZD�w���Z�Fg7������d�N�j:��0=z�����
g7��g7r������eH���DS(��5l�E���U�)����e�q������K���9Г�}~�����Y5�Bo6%��X��Ǘ C>��|�(�̱���TUEz:S�Y`$*V�(�X��z_� bW�K��\Zw}�/;٨�V6������e]%Ӳ�x��l.�����)<��І������<�6�=�>�z��笉�W��X�Պ:ch��ꑽ�횝���b;,��5����F��L�a�&"�Vz��q2��6�y�]zn~^���N貕�t��h�"h1�<��W�����`m"�]M�/����R!x�����'�U'�/^�H����}�'��~�,���N����ѩ���w�/��D��9��a��<��K���hS�i_v4���� s3���(腘��6��5��9�/��Ld3��t����a��a��l�s,�\`���%������%~�����TUU�g5F<��{�}Hi���+�@F՚�W=	Y}����%(�F%�$�F���ߗ�����^`}�{�����|̚Ǽj�(�XWn2m߰�0��5�.�.��u�U�w&��෴OߜV�`�tʻ'�e�S���Ҝ��q9=�cQ)��C�q��v���$�~(�K�q�kg�>|90s<ALF?�m�NR䚬��?�"�(��B���&��ƨ�o6[��G�P0,�e�6�tEzߴ�&@~ޙM�|s�=�D��h���Y���^�t8�b��ab��l�2��ţ��c�E����4򺎉&M8;C�.�E��D6^�������n�� �G?"v^���.+Ba�QZ�>�,� �W�Mv�����:��P�7�׉�3��漌.��ݽ�1a3>���}������{�d������S���r���=6A�3i��f��~Ղ��P����`m��1|{o�x��'+ʮ{�[>�4�3\*��-���i'&� ��*�z�<&Z�K�t�B;OK�x�4��m�U++{�J$�W[`�8�c�(h��$Ƚ+������Y�217o��YM���D�z	��M�*�r���ėo{ʦ�'� ѻ㴎�&(�����!��W�!ɳ=e�ؓ?q�b=�(���2j�A`������(��$���S�Ο:;�ǁ�6&�e �J�%�j#�`(c{�!Q��y���<l��p&S��h�&�oڋ?؋=�ON��y����csll��o�S��Y=��w���rc'�7�7Q�W����㒙S��W��K�L����`c���~"��l����6]�e������S���;���_��s>��O5����<e����?�׷J�W�5��
U#�g�˵�kꪵ_�K�[˄]>/��n~���)�]� ����W��F*]�L�aB�F o��>Ժ*�T��X��`��礊;Jleee/g1����-Ѯ.����Y@JW|HS]]]���a؅[fm䌒�N���aՆ7��U�1S$����]�Դ�$�v%� ��ǇsK�T>f�^�s��KRB��������R����=%� :��?���]�{bӘ�!z�n�=~% <U*)ruu��l=\��@ik�Q{h�&������1�4_����
� �cm_��g\L��T��8�lो)))�̦�O�t�m"���+.T��7��ir\+:��1X;�&�Q1�������q� ?��8���������ŷ����\~פ�!�Rk��3l�5��F����#��)��*���@��qeĬqkD�I~"���![+���
2���y�y��#��;�Z��O,,,���Q�u�S�!���S��'	&�}]�-��%o�����h�E!���q���lD:�*�l�?.]-h�Ф�!�IM]޽���v0��AA?�n�w�;]O�"u�&۟{hP�w�v,�6Ďj�̝���0�������O�=s��p���˗@�״�u�t�Lک����ħ�W�=|||P�?�ݰ2��Z���e"+���R3�x?���i"$9<�<�U�b�'�<�9�J3����Uݨ��S�dV�G�@U58��0�M�ՅD֎"<i�����b�Ȉ��4�5Sy3�F���g�'&--ͤ�E�P��|�eK��9��_�2+�W�'%�����s}FJ-�&&&^��s{X��&]{�K�ǃ���m�3�_���f^��9�P�d���s�D"#AYm�U���V�>G��Z��j�<�W��_���|1v���,���I�m9PpF{܏ZZa����o�?ȩ��gM(.;sP��0�������x�� \�y1��]��~��I��{j���Κ��2���K`�m��G����nZIi�s?W���(���z|KTA�\���=_���`�:		Iv�>�?��KN����\�ץ)�*jh�3+���ȥ����_~�i��8�s�{��f��~R����+�^�Q�l����Nڶ�!R�B�f'�����&wyy�u��J�4��4«3P�����Q�V���ӫ�����~��Q�N?xk�Vض']=�ai49%����o.��ݭ�-A*z��Z ��<�%R����Q@0Npm��_��?,x��.S�����(@EEXwӭ��츌�g�7�T�l���ƥ�Q��=�0EԄP�o	\O����b�(`r���_f���#a���R	�������GTx����.�nk��=^{��n���GY���sq������I?:�����G���{����������{=�����M����'�j���>�6g����蹡�S�5���Cc��g�����'E�ޢ�������O:�Q�7�}�}y
z�����̇ޔx��
�i�6�y��Z۠Uxf�*6bp��t4L֗f���ϢDGC�:!X��Pl^(:J ���#���/�ټlhh���h�|��o�0�.�Xc}}]�.�e
~��g��t8�����R���H\�R����;��t0���`��@�4#�PUE�xZ��y(3pU��nC"	###�]�����XT�Wk���G��Ơ�k��Dhbס��D{[[��d�dɍp^���R&B�u�K�q�]x�#"3ي�O��$|=�j0?�~i�2���+����kX�XSK!/�`�˜�m�s�}\	�>���p����[1Ź's���4�~������E�f�V�	\�t?E����>ań�g
@sىxL_�����{�� n(�Е�T�CQ�W���	���&U����S��uR?ʆ���~�����.�
��sU�������2��r$�e��P2L�V��?�$�:�B��;�S�Oļ�HŢ#<թ����r�r��[he���LH�G���#6&H쪂��5i��^����&#��9>����h�$�*������T�1�&rb4�x"�}	2�sQZ7F�B�S�7Ot������x��i�_~��A�[��Cl�L�k�*A����ԏ�~�(���V�?xz�P�ut\s#wqh�Ќ�j&�<��	��l�J
x&���V�p����T2��+���BqS��S�{�_��&a?p/��P�Ǟ�<L���$$�O�P��J\���@�C��&
׫Ȁ���x��v�ފ���;��c�8��U�⧆T��֐�����I�B����� �F��,h,h����8j�`�ۧ�4��>�nʌ�y
�.����`���f�a��
�
�X��c�勔n>���ܤ]��s��e�iw5�[���<�>��5h�$�̘�ܗ�E'�=�ocx�Ƥ�2������P�`<i
�hb�}�E�_0=�E����t �X�J����+������>_��3'�l8�u���o���u��<-]<�h\,313k����d9��-CA����g�����gʋ����:�����l�t�\�?��h��^�;7����_Z:�����0
]��/}�A�7�ũ?V���8���LĬA ��ly/�QR����*�'�o�|�{FO��� P��8��t4i��������/.���[���i���H�u�5j�T������(��z�(�sz�������iQ �(��Of�~x�Y�G�⨮��������GmZ���-hi	�,aRfA+כZGF�{:E3�i��$J�c��w����-���M��X��n������~%�r�N��1�Ewd��p���V�~�{���|�gsxN^�_��v~���w��:g�<I�����P�^PSk��d�MK����^�i5H�W��;N��iwe,46
�`g,��	sF��9�R�m�Q��Q��QOV��ե���a---��g���&�x�b�7�p��WII�Z�I�kO����D�����땆�!�R=A�h���D��� ���q99�	����C�/��#㛂�}W�D�����o����7���{��VU=���i�����I���26H����K(v��Ҿ��R�!��us�t�y޶�-�N�6���޲�<��3wq�v�rm�?<�3⒚���
5���)Z3-�<}/a�-UlR r#�7o�g0��U�c�PSss��'2��)����Ϟ�]��@'u]�~����SJ��}W�����92�LƩx34>��D���\�UqqqLӛ)�(0�,m�����cakpJ�G}6��N��tA�P��ȖX�?��]���M�853���-��NT5��1F�i���f��<Ơy����z#�W�C�ѻ���O�����y���f�gk���� Dj
�M�ZRv..�m,D�\J�����8@в��E��\A�c��SI�W;����&�NFCC���asiii\n.�_mp�%���d_l��و9�=
�� ��85�c��?�eê�B���Ka5���>�.�s��8�����6&�W9g���pe��2)Ϻ��<I��܁loo�[緙�4K,�A�'Ep,�KI� �hǩ�����+7����G����d.͟��5��O�v�P�P�0m���5�B��""����i2�����(�J�TɉsѼ�ȳ)(S����;�8�mn��@��(�wC&%-\nnnjZ���zj�C@�(���.�~����p>���6Z�b����Y������iKKK�{�������׽��o*���'�] =��0�]�ob��6<0 �r�Cn�),,�@U���3�1N��R1��6�8��0��1(������6���\RHS��N4��%P*�,�h�e@��3I{Ս���V�X�b���#�^z��K������n�ز�J=^'IX_��RN-����S��3j8����k��iɧ%	6o�h�؀�i�?�F��\&&8�	.�F���q-7�ԣ��%��Wy��3r�Z4�8�/�#ȴ�ʳǴ�������Kk���T�( Q�QE>��A�|���Z�	Ý7�i-�[#�B�=��i����{Qig]��¿�:X�ߣ����O�_�VZ�k*V3+?S~���y��C{��1���N��`�T�H���3�[��������@���Lq._�|�{����Ւ{l�l�ݞ����:����~E-����N����6��a����޻/*W���9y쭣���~h�ࡩ;=�Ю��g��W���:�}��?�>��1�,��S�R�����(�FAR��R��m%s�M�����N����P�re��Ocxڿ	ц(�i\Lܸr����'��e�ɇ�>�stmj�/�^<1��2�>�B)�zZI�Ɩ�U����Q�0L}Z+�'LY`~B�$��wm[3O��I�a�f6f��ã?Ttu���/M�'�����Zș��'�p�g8���W.�i�+�y^=�b�D���~ׇ;�]+��5�і&?p�ZL��M� $YJ�x��ŋ��<.�>k�p��9QS���]����"�#;t�I�In�dE�bT/�q��h����"�,<,�=f��QB%��2�%%���*W-���K�dJ����)�@�4��[+�� �^�Mr+��_�����r!��	�S��9�L-�󮻸�� %=�?,:!H�GCrZz=�����r�bU���W�і����gB�Ǉm�T+�kt�1�X�7ì<0�s�����yk�R�M`V��MQ�2�a���*v��8�-�l w6Ĭm/�ޑ< _�h�
����-������{;J)�xG,���;�0����|���~�XR��2�]hh�5>����~	����%�wV�����<he�l
Žt�RnoR��q������˸&�����.���(�;���f�Kd|[���sۚ�6�&�Mȸ�:�]����#�����0�V�ɨ����G�sv�࢖=1������>{#pQf#Tq/J�Efsۀv��}.�8����\�L�C8-x���sl�n��u��3E�rN�B�Bk�Vf��v�>��vx%�R��/�ha.}���-M�i�,vA�i���G��p�\6=�|)+��3J1�MmT���𢶅$� %:��j�������C��2́�!��%0�z^#R�"�R���}�W��-����ԵP�yc(�q���8�����,6�;��}��R;���n{�6�LL�l_���PO����cY��D���&���Io�8�v�N+#;�Fc&� q����Z��0�ѷKwZ�[w\��ֺO)��ػ��D���Z�j�$M���4�7��Ё�Dk;L�U��v���sW/TL\ŒD��1��na��@��	�a�E^]�cf�����Ą��o��ZkX�h�<�tj�q(�雚Z�ѣzlb#����"s_6	��g�h⁻ʨ|,ԯ���>Y����¹@�	�x�no4�{)�-�:1s����ЍYA����g'՗��5F_<�:3&99���U�VA!�	�ѱ���{|B�w�gV�m��tn@�7�ù��6c����+7�w&���m���mxIC��+w�|������r�im>�@韭7���H�7
�?n^t��]JƄ𕃚�/��IJy||<�&�QM�з`=�l$�|�!�v�[���`ͮz��9��x�{�ill����u�(4�#�Zo��˃k��G�J��[�^-��R���α�J������3a�@�0d��~��_UKt��~e����W��b�w�5��[��l�uQ�猱dN��>{_����\��V����_I��t�pׁ����1��tu��jR*w$Hz��|"��rɉ2�թ
c�&�>H$~f���3��J�暏l�U��z���_��Դ@%4����1nݵhJ��7�u\�]��!��vZKINvO��`����a�������A�jod��K�h���t�A;5qqȵ��/�� �Q��D��|P>b���YONr��5wM��a�3���2����5m�|�CK�v���I����>E�ѿd)0K#�����$��b�l�+�Ƴ�s�Ό�KmP�7�F�W4�S��#+��U�ۓ���b�_<ǁ�B�qˮL��ƍҦ�6g�D춓F)[I�5������j_��\7'�-L�,�˩z\{���(4L&d��F �N/u�7윢��](f�*�c��W�5]��;�l�O[�t��1Bh�R���m�da�^�\�� �������r���cն8��RJ�Ȱ� =��\ ��^��Z���HM�������>�VG����ܖ�(RL(>�"��	K���b&���"w�љ/?�~{��.����S�;/G R��&�W{HG)D�	?bxtߪX#��z�l�2ޢ+�Uj�ϙ��1A ��gw`�="}�� !񽍁IZ7j�l�>�*D	g��	���ڱT�^IV�R(�W�H�b��:I�4�}�x�\���ꚍ�~�eϙ�L1�num5^F>������3��uɱ�2�޻��R�W	7�9�OZ ��yC�5|���w���`IC����XV����<���]���q*qM���Ę���p� 0$�?]S�����X�أ�(,E���]r���%�Q��r�%}T\$^]\��`$j�Ї�ߞh��!*�����!!��)|F��c>{�[��他8��*���0��/I>N�0Rb9�g��V���v`k���:V�VC:ʖi��B��%��>r�,�5�[�7i*Y�k)X"W���߳'<+�p;*�*�6�W� ���u -~�׆�RjP�;E�&�k6wU@�Ss��#��`ЮCc��;X-5����&�0BB��g�S��C{	������c��{%~�
S�!Y1Lh�!���
��fx�{CB�̰u��̵��[ޮ�,K2U$�����;�O���b��x����G��%k�8�������y�D�����.����gQ��S����3be<N���uxt0��Y��&�Zc�j&�vC?ڙ͆a�@���p��|�����`?�+�0o�``�a糀;�,�⊢�sd�W��F�5�@�%+�=���.G�S՚vO��X��˫5:���у���X�����#�+�S��L��B_ɗޒ;�gn���ڀ��a�`�!��iږ��L)�=����ޡ��TN-j��5{;�C��k���ǸB�C����3p�"�0�R�Ƽm�jձ�ݫ�}̽�ްf��Y9�N�.E��mX6�C�g#�]��7�݄|�bܟ��g���A�$��p�u=���@�W�.�,$,,,Y�[��i+2��G�~��I ���n�w�\��Zn %O���G�)-���$J����� 't���ٜ[q㙅|�پv�J��������,#����7����d��_�_�����+�U�k�P�Hi��^�T��i/���7{�.��G��L{��1�k����s0F�1P������L_�7�����c�l�(�!�Ѭ�/���A.����\f+��ॸ����l6@��!�l{K�1�?17w�?G"���@�O��|��	�S��,�-����͝9s&�ica.��t���w��F�J~}|+
�˧~��U_t=�k�6���@�$t�ڊ�D�`����}+Y�;1�D���e�+t��q��?�s�'��j�hk:��2\�l��z��^�%/ݶ��C�3����ZBU��]/�h��X��R�՞λ�ܿ(���nىbly��IrB�4bi=���b��ٜ��������1��a�{{�6�c�銱��j� �9[�2�HD�q��I�lg�bq]���"�>�1yG�]�����ֱ�!}�W͟�]�\p]�qe&�є�oJ�Ɨ6b~�{Y��L���"�bQh"r��@r�a �d:�%a��'FY�YEB5#�JK�?�7"���6�Uʅevf��Q��<gm}������Ɔ�#ȿ����;=\!�Aa�����9�9(��F�`�3;�\Cn���ηr �)�JY��
f{H��T�@���e�:Z��[ޟ��|���3�C� �I6fu�+C��w�t�E ����]@eK�
�[�@�e�<����cd7FYcع����*nXG
�f�M��
��؉L�kC\S�e��G3��>7�&-x�lXD�7�Q@#j�E�C���
J��j뮇����V�ܬڑ�����j��pp���;�A����ݼ']��Jn-;��A��E64�NR���.�������mv�ܦ��3M�tc����H�x�?o�QG���@�3q4ut
��$}��C��/������LlV�Ǎ����~����W�#��e)l�]�I�Y ���
�$���	���"<�`>%|��Q�P���66���5��P�H�Z-ƠR����ӹ<�����%-��r�>�4���}A*<��o�\�,����N:&M�	��䗓L�JR#���a�@��@�';Mv��ԭ�c"��j���PM��/Ta�;��ɺ��D.��jxɦg\i��+Q-���~��&´��@��T��q#�1].ɓ�&E�@�w!�$/D�Ƭ�Юs絘��d�ԇΥ����r�!/��ݽf���f,�d�/t7��y����O,���V��Qu��KJN��>=�;WWW]�F��t1~U��g_ݤk����ok�G"���n6���_��*�Z�$]�Zb&��ݶ[n迯�k�=6�|z�յ��Ȟ����_�R��P1v���y��.��e�p��-Ǆ�J[Su���S|Ձ�i�v���+�������e{rE�(
�M��wT7�&��R�b\+��MÆ�7�G�"u��L��M�$�����K�R88��s�D���";�F�D?���o�{�
�|���/�|X���
u��-���>OĵU>�}����� K�;���@(EM���7M�uԋ��=-N�����T~�
��9��:��`L-Z.-<���ɶ��j0��(~\4���|�h^�����v��!�jQTB���r����
�'�L}��{bpf�.i�j�X)^���	%�/��p��)�f5���o���L�Y2�	����<..��^���S�}��B�纳vMm���J�����ؿ�N�@�[=�2,���%5�߿T f�%i8տ��ޏ���!v7BŪ)�>W0�f+�P�!��$'���i葓>Oq�����
�q�i�e�����͝r�ُ}?���f�_p���#�r��v��, ��p�&,6�l\u@����9@B���!�!��-)-ݩ�4���	Hw(�1BZ��������W��?{�m��<�9�3�$ˁ�d��f�bS��2��99�Ǒ7V�Ő⠠ Ú�6�瓁�J��ώ+�B���Ty|�,����zAk<��`��Q?�ԶGgnz!�Ly��G�r�H�!�6� }��y���a/h$���鈛�Պу��]3�.��+��y��p��ן�Y�=�R��-�&�^��wE�R	�l����t�R��Br!����F�|� 1>�ߴ��:l���"���İH���cDvt�  $(Ȏ\q�k�{QM��olMl}�#�3_'<A���)���?xA���/_"=���������A�b��K�v]⩭�><�����o�^><q�\�M)���s����ދ,�<�)�Z	ۛ�������E�{��i,����Jd�Y�6^$W�@���l3�em�6��=�>R!�I�Pˍ��II-�==�͎ۨ��8}�RF�*�k��I�Gh\���2�R�E5�Q�E�r�L��:�<��3+߸�UZ�ha�+L�\��|��.G���0�&4H�4쩒����6�~��ģ���.p�2dddd�������n�W>�P=�V�1���=FG��=�G �,�<�^��fZ����zg����7������<L �z���˽n��ۨ{S�&`��� �\wW�	I��0q�h��dn��L�b�z�����&1�֪iXT����y ���ô)<� PmGT���Xq��j�9�Z�XIk�|;��:�WU9H:�b�uջ��"��U�Us]o��a��3o*��lޓ�v<�R�u����50F-�{B��*t��u�uxc?�2.��<���K��Z!|���W6��&�8[=�k�)7�|u�9'���)���m�)�!j��[��d�4���>B�N�%�z"�	5X��E��)�
D��i���ȃG��*�YTמ�Y��?�~&�́�hg�{��K[�_��$�10�^�*1l��%��e�"�("k�%T�x�b����RpRg=����do�|�)�\W~*Ӷ-+�����b<���/6	%01���(�^�2�9��[�~�(���DLv�`�^ {�������o-��5/�+��HH4�֙�ޫ����;�����Ω0�q�.Q��	�#o�-�ڀ
Hz	7͔i���z�s[�&ϫ;�O�����������5CÉ��Lpu��R��8nC�K�b���m̥��w7����xf03~�f	�S*Yϐ��E`�Ges����nr�@��.�Di����sԣ���R࿟=կ���i;J�Xv�E!d	�C�,�k
S�#e����$8��ҟ<���v�h����`u�#7��B����?�D �nZ��˗tO�3)WSk��*h�r��~~�`\�èm�+}l��?j�=����5p����ü�HP[I�������Ti���pFz���M/���w)0�6X��6�}����J^ޭך^����)-F��n�d�lY�gZ.��(�	,��Au�]-�i��V ��.��g���$�JmC�{s�c	jv�e��-{��狝��R����-oxQ�?��I�W�J�gֈ��h>�#�d�a5]{��h��Hq�WJ���=��Z*˵Ý����U�[�|	�p�U��q����dypB$_�lW�~�`w�y@�Ǌ��S�� 2� �H�����q�J��4�������Oǘ�C|� ������fr�&�_{��!��R�cK����N�wXEa��F&w��G��5<���(��pO[Q��)�Ә*��J#w?�t�!@��n��������-�Y�\ ͘�f��>e)�T�8�Z�L�.��p�����:�^I��N�kr�S���R"�;�D<<m|�O���]�Ƕ��򈛛��;�1�0���{d����^�*��o�N� ��Q�h�b��zg���<��,)-�xt���?�
�-��ߖ3���O���O��MV(�_f��&��{b2�چ>�]������|�^:@���Y��+�Ѩ��@ъI� ��$���=y�9��$��B�:�V;�a�S~�Vt��m���}OaAa�*s��uo�ρm:�c��Z�{Ϲ��vێ��6D����e�dLXC��;e����+F�扗�ǔS�7�'������n�^�\��)��@�=����UR0��<�X��e%��UU���*�BO�m�Z��N�g�~�z���eϢy�Jk)j��t\_�7��ͧFz����Q&т��\�U�e����BG�ߴ���%��˺�X��eR�4g�x��.�&H��(󣞩i�7�J`�.\f�S���ȇ �{����'����M�qѐT��'�[���ޒ�Kg9c4�!m�<��Z����B��Į>��	)����b���3�cnZp��>y��`,Z4���M^�ɺ���J���+ύ��
�hXj��l3�q�Ԯ��$$���b�{H�?�c֙��^R�]M�).+709,!��0�xy�C�+uۥ�_O<�&4�<b���;(�ap*�n�"�s!��^�Ek^�%�Cx���QS1D�z^3�OB�Ӈ.+�?-PiN"���?���X�v<���E�?S%%�_s��J�Gx|�,�@��}Ә��	�s��}LoqGU���������7�~��Q!7�Ã6�hݎG"�_�ݠ+ s���Rc;sI�<�n�3!��F�F���6J�3h���RQ��V�(K�A��X!Xx��ϧ�.k�J'6m����f>�EY,�8:��K7�r�F�w
�B,y�*�<BL묯�Á�%�^u������5�j��$��vf]<��.=��b���l�.��t��b��_�*s�sp�h]Jb r-��[�)A����U�����*�T&v��Jhn�o�e"��tU�cA�Q�N�g�*�ݜ�0U�9��WFs" |w���̶����a�bn�Yk9D\�@��e�\)!�p�tf�������5�[:P,(���37�f����`�GN'iդBGG��<�F�un�E!��f.ϓ0`�͏ȟۀU�gt�?�z��!x~��Vu�Y!��~@���<1�����MAǧ�l�:Ky�0˗ �9lO��67-�P8�G����n�S	�54������QM"��Y�]�sυ���z3�� ��U�����V�r��⦡�A�B�D4�߲�0�����IV_�9�*H��xW�B�l�d��i1���0zw�{,��+�0R��;�W�0��O���lm�
*1�B,~�K�|����-�l�TZt�i�W�i����R���t�[���FS�nՖ�q�xx;)͗���D\�tUl����Y��� ���œ ������DoT������Mk6�T�Avr��Bc��vŮ�1�'���.4T��m{뮇bi�u
��/��V�����>YS]�廊~bs��{�YF?B0��ER�ظ�����dB��pc��`��j�tenm�L	�H�_��m��323��𱕿�K�}��"0����WU*))�6�D{0��zII�PJ;�un��d�P&jj��7"�0��n�/��N	�U��|o��_�D�i���9q����n3��9L���CS�v���8
S�3}�<�*�kʐ�S��l��,�ŏ�!��w�����@Z�9r�v���V�8���>�n�T	8@���4���6hzD��¯��<7d�\g�Yj5�ӗ���k�'��RAZ\�i���(wr{�ӗ˨�iN�^��5X��,qr�:�Hy�4����㠭<��-+�O,�kz�XsJ�,�vz��SF	sUsH5�%==!��X�������1��D��|&������v���r�Pϯ��|4��Y^����kҷ�7�g��7���W5=��A?�e�vL �dYuzZZ�*/��ottb�����&]�D�ؿ�b��썴��r�q��7P��GS!�!e-���6	��+@�����{��0y�"�AX���k��v!`DEiTb^����Ez�3�g���Au������y�Ҁ�W*�ގ�z�/�_���@�kpC���+a޶��w��s��k-#�� ���
L|�H�������]ܸM��bo��d����
�O�h�t�I�b�;���\���{^�i��[�j�ey����)���
����au���,�(�A�y|\��j7'�u�C\��v��j8�--W�<LNX*VD���:\��(t�e{��jijR���1�1�"őa�q�k��[dPZ�W�%.yz��7`;O�ܼ0�������R��ٖ��b׻U�J�zYf�hau+L���EZ�J�0�#U3l���Bn�h1����.�r�R�:���O���Gݟ	�����A�t5A�8O.��І�8��6�^a��v�i��==�z���5�nx��@rNV��Cc�S��|:����^h)f�ot��.Xm���p�̅��F]���U���1�Vy�=b<�i]<1Y�R<Y�b�nk��X;j�мء����&��fM�E�%�=7e{3>}�����&����wb��Y�[���溦r�k���&o�'?����1C�s�	y�O2
�� bX�oO�9�b��׷��w�n����p�C��]�t-�u�s������(���%s�<{�g�R=�ݭ�*�Ճ�"�������-w�I��Z}�Z�tp�3�~�Ӛg�7b�>���r��K�J��%5�ո����8�K��,x�.n��6��Zp.�/�˓S�����Z��6s�A�-�?�_��U���j!�@�c-0&k�<�O"SZR6�Z0Oڡ��?.c���̛��2b�T��x��#��f�h�K���3M����E��a��R��yP��+����+����������\�8n�ê�r���+�����%�tj���~�����������٭���-Mi���%0�(�ђ�l�RE�HN��:���g
�O5�nH{���;��By�/����.�����,��e�wW��	ɬ'n���6֘�Vr���@�O��d���"R�:{e[z��S$��Lȴ�m����1�[cY9؍n>
�$�����>��[�$��s[7�w�{����,��i5�w1<`����v��.9JW\*Pd5<�f�D|@<{39ꐧ�i��� Z��hCX�O�M��fk9ű�|2������t��I������T��XŮ���P�B��	�J)7*fS��I��2g빥YEM,_�ֱ�*6m(}�s��g?s6���>��޴\9�K��:�:���c��g2]��"�:#d~�7�XYٻ7� 53�Ͳ��N��/X��>��!
xRo:8;i�Z�5V��w�J�}�o��b�b~���ɓ����.�3݌�")��=.��� f�m���/�a�w��*�Z��[��g*ىf� ��4���K��멫F4G�����O�v�O�X1�(�g�F��E��$j"��p����s�*��-kM�7F�V���J��\zW�\�d��6$�b�����>�(�MΩ�|�5n�ԧ��I��K��c�]��s�����0������?e\�h7�c�E*?�PE)�nji�����Y*U=����z����V?����pL���R��M�C.����M�ܧ����ΕP�i�T�us0A>Fm���c�6��.���11�[����w9����;�{F.����g�V���/)�%��.� ������WSݲR;w�)n�1�-�?b�����,hgiq�c�J�2k����X&������Xm3G�ʻ����{
�V�_�mV����#FS@p�h�=�����AD ��wj�ANyݸ�x+��ܲ�h���-KL3��n�M*�`޷ ��ﴢE0 ��V���zøX:�_n�R�#	�ݼ�6Q�%��a�O%��>��-��E���iEj��$ߒ��c�e�6�e�Qg4�5���d޳P�jܡj}��%�\m�A��.���9GGKy�-�qah�U�Opj;ͪ6�����E��2i�I���2V*��[3Z������I�轸�%
������ @�q�WfKT��V�Q	�����2�^��w<n���{*��-�v���_鎉r_)���\�ɟ�W���L�)�8�a�3�@��3Vn�ji�^^,Yr+e��' 6�/�4���n�;�w�8���3�#��b�Gm�3������u��#!��Xt�U����XQC ö"�,~��u���+Q��'o��{kOe�h�ŉ�������|D�L�)���!�b�>C���n\��8
��һ@��a�4y�q�kͶv�jV����X����L�aTk�C�L���.˾P��X������,k���B���}S���������
QTT��Z9%%r44G�7�WMt��Ϟ�;t��a|���h胸�N-}Z��޷}ު�)��/[u8���Gk�O��?��(+S�d.J�IZ�|y�-��q1^F�E/���Ϗ�oy��c��p������T���@��+o��{�>��{.%�y�'rT������}��>���H0� �ݫE��m�|��qV,
-�8�c~2�Q�XQL�Vz��.s���������.�V��n�W�{��M5�L��2'j�:U�"uD���rs�L{.�L8G��c�����u���K&3����YۺA�09�Z����������0ѓ�$��/��'�]���9<�V�Ew�DQ3NV�P���53��CU��ӳ
�ߜ��v��qnc���'��k�����Fl�+�#�\63���f�|��>畵2Ss)�d��2#���ʤB�Y���^<Ǽk����V��K���@⻛,�^Vk�H	�~�����K���,#|�`��5�o���>�Ғm{�B�4'�l#� ю����B8��� �pjk���r�<!x%9^�K�I�g�z6��#b��tQ"U����V�C.T��(]
�-'�ђ�I�Ut���H�YJdL����]���Jz,"m*���9hR�>���}�Y����c���T��0S��ဩv�OI��g����?v!�b|��*)��A�B��b8��S��[�N�����{��ՀF
���`���A�j%d ��l���'�̀Ϟ�Y��mB U9���0^�G��+g�����~�8��ü������d^�񓾻�&�#�r���&��L�ni��� ���藕E�[�6�WR^2���ϑ}����!��ָ)�\88�R���s'��gث�O[y.�c�M��f��X�%�Wj�/g��v�7[̷{���+�������Ëk�d`�	w@x[WAt�p�k���:)'/5i�0���iZ1_�*�i���b&�&���.�}4��;t:ي/ l��퉋Ǝ#ŝ��(� ��NkhQ�TϨV��D�J!��D��&!�����"fcS�2���ɩ�V���n�x_H�զf��-z���[���L�0T,[DT�`�$u4����!C�l�Om�(���9��^����k���
3�!bz���)=���<h�i�n-��q��uHK_�;�ƴ�_%F�y������4��j��u�.�7FA��iߎKXٯ3�T��0f��j�d^�oQ�@۞9����:U��Ė�����\*@���\����)Mv\�1���:��d���JJ��gu-�-��bZ���]]�<�Bc�0�ˌnU���7;�)��eo�a��A��J��}6�xSN-ejIF1HG+.�ŋ�긊���*
V$*`c�xz����1��s
���?v ��w0WG���]L���}��4loM�?�0�g��r�!°����ARz�AO��U����k�D*�����Bt3h�#�%�nU:�gB���'��,\�6��b]��~��JnvK!Y����p q�����O��	g�1�V�[?�G�qS�ZnOT��x~��2?����_Z�up�'��M#"w�:��PFH�$z����Y��w�a�b�]���U�F,�z�c<��!c�~t��q|U5�o���I���}��0@��"㪹�+N��w�k��2��$(��X�y��OW-Ō%Tq��������9���y�j,k�\=�a-�*�����`���7_�8>~a�g;7!��C�hÄ��N��	�����G�<zGN�:�f�.
>���< M]�W�署���,����ۧ�Z\��Ԉ�R5���''5�F�R�>v������I�����zU�e�$��Y����,��R���+1fRu������֤�/���d�)I��gn�$��#>�V���^��E�Gx&��M<4ST{��ߥ�
�Y�3W#�汝yG���c;4�p�"�&��aa,�H�k�U%���Zm�w��`�v%z.�}��^_�KR��o��	@B�
��`�����|�+��)flL�� Z�k�F0	�H�Q#��̣�99M�䷾����.!$$��<��]3?~��������cTB^��SS��m�g��-�\��2|�T�Ղئ�n�B?�kDœ�Ê���o���j��oج��� �
J}��γc�Z���{���QkNg��L�f���y�W�ߊ���'p���/�AroS��YHȎ8�PІ3��9��|i��oIr�(qHH�� ���2����J]��yL^H=�KO �Kk߄l���ۘ���V��~$�`F�ܥq�r��Og>�y�����������#4���=�ׇ�j��_�I=�`�]j&�k���b����~�G�+��p�Z�Q;Qy��J��{�~`t"իd�XfͿҩ7-������gB+�Y�O��?�# ��T�/����E�h�L����\�T`O��p��T��ڜ{�N0
p瞧��ޛ�������W�F����km-�m��z>�������!2g��k�[�6+�ۙ��u����?	4�}����m��CKT���B��'"xމ9���]=�M�G��y�ĥ�n��\=�3p��H�+~�g��ʍ��/��9@�K��+��C�#I�'���w�Ͻ%��XJ�"A)���O&<#6w�0X$ar�Mh{G��M���lY^q�9��)�a�M�#K�J���5++;�<`YcG��dq���V�~7��n�'��|r��b�����s�X���}����&)�Th�OW� !mU����eA������a3y�q3�r��GNmO��h��R�w�Q�G����ܨ�-����ՌE�fX��`�0\�C�7K���:D��8�1��a�ϑ���+����^=_Ǳ��f��3ՎT7��*g�p��{�F[,��75�I?[ޅ�s�"�@Ǥ��م����Lܜ8������oٮw;j$�)"Y�/��E���<(�x���%��u�_�Y�b@�����'���/�ضc��0��<��XUX�I�s>g���mOn��gWX�1v�42<ܙf��kL�@�����%$�HJH?77/�1$�l}���.���f����9�cQԶ�wq'H�� �����}��E����Y�Q�4A�x��?�H�щ��D��t!5��Gc�V�6↙Zi���$�iȑTy�	��u�{��XsYa(�įq�&���<���F8ڛ
_���M`1B���ƀ	`�*��j��*8>�+�" 1��ˆN�*'� m�t_�Kz�t��X�U�H�e�ԊB1���k�����%��[�53�|�6���v6����@ �7�r�m �	J��6�j����$Nc=Zԝ��Pޥ�!�b�������|is���.ڢ����Z�G��2`7H�Y�2�%0��H)���jN�eUh��
~Ft9�u�g�w �ӎ=�
� মS�p�Y�Ϧ�ڸ�ѣ��������S�E�te ���Y���5����.�:ʇo@��i�b;e�]�\j;z�q�q���͵��ˈ.���cF�Snn���<q��m���oM0��ν<x�y����]o\��
o�;p��햡�D�ex?���e��] ��v���EJ`��{��w9I���R## ���-=��80���
c̬F��&�p�m�'��(1�g���R^֠���*�F&x�e���NO'�kԶǋK7��.�`��1=�G�R�][�s�J����%|
$Y&�50�G���\XPY_���������q�qU^��/�$1`�^ތR���R��q��3[ �%��k�ߛ�~�Ȏ��Q����($eZ#q�JY�~�� ��!@�A6�]�J��p��2=%bJ���s�kѵYRw�ƛcF��12|Wk 6�8��.�s�Yo�iR>�
���7mhxPl�hADBc-��<�@I�wQ�J��y�Nq�t������q5����1��nx�C��\�nm�MC7��J��<�b��0���9EYII(,��_�F�@X�P�Vt;�2[�lh�a�E�̉[��~5��G���]8��1���Jj {�-E�^��]�Mj��A��&=�n�:P�6j��#��:7I����cl�g$�~����Q0$�^�NZ�撐P�2=M/�r쨡e��5����T1�d��a��6���h��-��Rk+%�Ch��$M#m=MN�vS*�������Y�]��%��!�ޠbJ������<Rݸ�����2�$��22��L���D �-�,��r�'?����y�a8{��*�P �A>���0��T�L좄8oa��	��N���AP�2x#*�ᶔZ2t
o�+�m@�|�Mд&C��_.t�౏���{�ȃ���(0nu��#����᧓�ҶV^m��>8���f��9i1(��P�@� ��a�װ,�gW�J��6�z9�?V��x��o���0�Y�bk��>�J�a�3ȫ-,���x*��8kĂ��ñ�����<���&�ɘ¬�~�&���*���
��Y�Q�cz����O>�w�냿o�mFD�����Eek~�|�$��p�)��)	��Z���]�Ղ����lM�.��B�n���W��+��N�Ę�~���9 i'ð��v�?x(Ml�l^�+�;�S�4QR�Rv�eV��P� ���06�WI�c�u/�-�^��V��fj
�fpoʫ�6���-9}Z�8,R��\z�������Z���o�S�}ԓ��>:�4g�g���\υ����� d/<�/�N�L�	H܆�������m�5M�ٔퟯu7�-�RZȝ�b��ŭZ v�8u�~��ƛ���������g͍! v��@�?��_���G�lf���=�2J�t��38Wf	�k���U���ފ�.@�v̖�qA�����J��'����u-������Έ��1���� 5���ܙU)D�收�0�8�#<���=8Q��8F��衙lx=?�ew9#��?Q����YO�;\]���j�l&eן��r����We�o=R_vQ�׆�+��W}ve1o�m��u}�f�V�N�q�^6%�U��0"l�2P����@�V�uœ�<Դ�/� Hg��нm]�5���[��gw�]a���k+f���C򾔼WBl �u���6��B]��Q����|�@ps߁&5��l1��_���\O�$��9��&Y��٩�|���T��H�@�`���T93�B4v��^���f�	ϗ�M9XETP��yCW
��6����2��)�y5��
!6��4{ {�3x��VLYĿ�TBSD6��P���=�F���ň���0Ȍ��;S��k���f$���F�%auo$�2/g�0_E�8X/ϭ���.��o���#8Tj�W��H�f�*^g|)�� ޝ	\"(
f�yrp8;��=JV��)�����7��{~�c=ZZ&V'n&_h����;̛������pD�,U^���ĉŭ�&ȫ�����j&=}�R�Ƃv��r�����$��K+�De��'m�ӫ�_��P1L�9�qwZ�e
9�<�k�n7��v<�n"�l^�+��#�A����/�i'���u���L���5�w|l�5~�c���x	q�O��s���&�Ćz���}l�`�I!�~���A�h�D2aƷ�b���q|��%����;"�8�,�j����~G�60+����4\�G�9h��!y�9u�5�OJ���_V�L�W<ef��+hߕZ8j>�YE�g�3a��T�MY��<�#�6�I^���Y���|���X{�5A&��W�>r��ݔ���/�;���C=���lZj��f����\���������K��HvH`Uy�H3�2.6��8��x��
&<�N!�~5'��WEWb����ZK�&C�=��#�or�UU��6�Y3�>��K֏���2�-�{/��%����i��#m$��V�)ec���i�ѻ"�ޗz��꿖��iVݤ�7z$�;�l�ҭ�h@U�W||�$�+Z+�ҜRМ�7���R�����Mz�X���팥8�x�Teni=��~<^y1g���s.w�y���c���-,���S�E���a�i1�<���S��-�����4
�1M�!��۵^�x�Ȧ0�N)}"�_\jv20vW�@�ԡ	?�Ŝs��EOI/>����L����|�ao__ns�^�����2�sCɉ5,�P����"�O�&dX'�V��M���jbu��W�3<����y�L��?I�;7���	"����Hw}�k7�����4���)ҙ21)z������|<x�d^�t i��%��͙d��"&����08J�W\9Kf�]Y����M��^}���1�R�n�U/�Q�)�c�nr�ӣJ��\����jp��t��&S�FQ���}1-/���e�lfVn�A�V�C��wVN����Un4C�X�vò�e�ƶş>�p�cbbB'"*MvE�~=��%8!��|�7�A�ª��K��C��}��bt��D�$��r ��Hf(��j��m�6�]���va���O�P�2		�b5��6o��$����c��d�φ�o�m�	Ͷ��!2~��H<��u��v@@���"6�eV�Ʋ~�ͽYd�2�b�v���p�e�Ì<�fvs�J��^��dǚs����,���ʄ�/��?�� 9����'M��T�� w)La��}��2��_e�F)�hl�PF�����,�H��A^A��p��h�߳$k'��T��`��T��A��]�3C�W�~��D��F�ʭꮼ�0/8�v���T�
?������+�[�ћ����m[�e`�z�;|�]�)5�n����s�SJ�K�χ�k�t�8��E؉f��B��#��n&�nhڈ^�4ˇ����l�r��Z��u���%N�E�&E	���`+��w�ݞ1��k&��&?i�v����B��>���*ZY`���7�Fo�3k.O���|�����?�+bK�����ё�&�:�u��]jm�ƷgcӼ��C.�f#(	�s �����)��H�N��l	8��������۞k��x�wkA�ڽ�{}�7��n�3։�Ke��f��:��@�!�/���l������X��D��h3] kw-�d7D���Zd�pk�_��mJc�ʱ/9��e��}}}Q��(��m��Դ���9�� �T1�&����5Я9�}�rV��L���i��%���I74RaL��S�TrQ�v$�G{�` ���l9o�ډ[F#�*��M
0v`uX�E ������8T,��Ce�@4NQS����Ӄ�̰��û�K����*wf6�5�Z�(���a���>�L�=����A�q��M6ߎ�ǌ������	�9���V�8��/؛X�a����ðae�G|��+�\��+i.J�����v�4��ld��z�l��&��UW�	o�a��v���0�v:w{K���:r�y8�$gټ�~j�_����;�J�we�K�p
�_�v5�?���K��:�����}��]ծ�����_R.5�������ut�Rt�ϟ?��@��[>�U)��D&wjg����x/�@>}�J~1J����aJ>{*��U�h?�`X��1
��`��+�7~�tNju����j	�[��܍���©�r$��R�b���'u
�no��J�>IZ�=_�J��2��B�s�]
?]l�����0�������7_�Bg0y��_���ީpw�
jP��uG&ۛ^�r��=pt�� Do�7k�Q�J$�T@kE�i�Z����M�Z�~M��̋)��e��ؒ�C&m�N��of��A�TE�_���|n�����Tq�>s7NY6�t�-t�Γ.������N�j�d�5�o�N�Jz����J�Y�s��o�̃h4C�`���F������r%v�y:}��X2Ia�˫K汏��ff}�$�9fCi�a?�ۤV��_T�����
�S|gv�o�35��N鋉��7G;3�?]��	��D���"�̚*.��\�׺���;0ǫ���x�+m�D����W7���������:]L��ŏ0����]�v��A��0�}8/��@9\-�x;~��g)i^�A�������R�^@��{��'�������?��(q1�5̈́<OK��_����O�h��_�����4�ikB�ۻyll���	��(��lk�8\[K+)�a�������f� 9n	R=�L�0W��#�= �������ʥo���su�����)������Z>p�U�S+�I�4���?���V�B�bͯ�$S�KD!��50P�o�ܸQ�c�	 ���,C�'�͎n���V�~B�'#rwj-�խ�6�$1|��X��R1ػ�|��2(�sAAdr��+TL0J�
��1�ҩ�n�&ڷ�O�s����[���s}|V_�7�*7��6��Y��x�za4�9��:�����z��oL��$����p���`��FY�Pj�yo�^:�.j����˻~�~�3�H�d��T�,�D��`��ce�iH�����U4Ż����:~/Ȍ��h԰4�l�hu��wl�BZ��]����!)��V�$R6{^~:?K�4�	�p�	���T*#'G$��@rD���[N$}��\|o��uRp��[Ae%%|���c�#�x^vş��kQ� e�m䶷�Kxz6�}E��_�<��o�9ڿ${�ZV_���!�74Ľ��^i��S��j����#�Aq|n�
}&�B��9k���ZsÎ7]�j�����.q�0�t���[���?_�]x�=���?O� �N��].�긝�&J��t�;;'R���������� I$C�4E��I]f����?{PA 66�r�)fp;p�;6&f7�^#�����4?���z�4rjkk�8Ɔ���5I��ٜj �� `�r���iE�y�p J��Y
�p��
U�j��;�[bl��(���X��L�g���U�� H���**1����������_��P�j[qUW�0~�K����3�
F�+灡�q���}(
����-�˹K����]�<�%D�f��0R�#�2��B�� 1:"�ٓ���ŉ)�?G���㐕�(�g���m�������;ndʊ}NDOM-/Y����0�]eG��|!�pְ�LK����m��BKK{���A�3��篦b�܂��
�]����W}���n���n���сyi0����o�!������N���Z�*121��8q4����q��Y�e���i�V@UUU�� �L'�"���r��:�PN���ae@FLL��;�]���LWm�$'J�#����ģ��d���Y7�Km���5��_٨i (��%`�B����ɤP�T�n
�X�Σߵ��1:����B�����A]���m���%�o�7
�=ޞ�������=�)������/ �#&.n;���\Y8!���BN��	x�؎"C22�ɗ(����l]�}�l�&�m =T��TJqy�q��_3�����Mٓ��o.��eJ�Q�d��{*��l)��{�XH"Lb�1�1,�c�����o�ʃ�DE�2wL�� >| i	T���.����%`��o�HO�8{Of~G^�VMK�����à۸-q����;C��?��Af�����:_�/��c?���5�ى,�G�!�lڅ�tRl1�
�CHE��$�Oң��v\i�}�.����)M7��a�H}T�:��۬�s�%y}� ��1����~	=�L436>ceWz����i
q���y��SY��� !)9"K�������S���%������%�O&aP�ҤI�ۢ=�B[@��B��Df���]���<Ѿ��gg�ϧ�!����Y;0?>��P�O(����	�3ɕl0uD��1���~�s�ۡ�ah�%ٛ2�v���{8�	Ƀ����EEत$�Ң��q�q�'m�MJ�q
����i����G~((��T���B��?[ރ�L�M>�~.��±洬l���$,����ӌ��8�βY]����d(��=?$,��8�l�K���)�?'c���QoF:f��F����`��~'��J� ݹ���ւ�̴B�A���Xt�kY�l��M.��E��*?ĹNiʊ�O��c�w�ҿ�<�t�(�%a�M��!��+{A鲴���c�t�1�(��͓O��X$zAII\pppd0��J�E�h�,e$���j;�#�L�8��j�d�
�T)��9Z�; ��zb$IO�#'M4����7f�s�)�۾'�+������d1��@D�=��J��D}��a�C�/ O�F/�ݴ�-����WSL|��s�&!!xc�D�9�����sr����?�,�14��\s׊�E�_g �� �,���V�ȟ�����<�$��YJJS�`�Q'��	���T�[��}��io�΃�P2b|ĳr�K���Q%��P1�3g'�{2d5�zj�YRJ��f�sN���Dt�yC�����m^��?�v&m ��N�֣eB���D�wL��һ�9D���#vf�f�de�:(���$s�aTˍ�H�#�Ic�wr��W|$=�y�@Q2��d|!����������}��݁�� 9����"�"�j��|pD�څbPn<�6x�f{&��D3��(7�ȸ�ԏaE���������ڤ ��n+a��q�h�Τ�<i.[b����)Ʈx�����VAq���R�J�w� ��4�/-�����нXxm�������û��1��{�'�R��jj����C�����j{[އ�RJ�������!8��Zܡ�
E
ww/P�wnł���o��{���/��X�df�<�<3�w�+��&���a)�����YO2k��p��?6���`Т��lH!)�����VnYʜQ��*tP���������%:����NS8O{$��Ƽ-H����c��������*N	�螸Ra� <�c����x���=�����{u��W��MD�g\���	Dhn�u�)ַ�ŉ	�Toog5���d�}�����eag��-k�N�?\{�t@�����4y�z ��x��l��k��1��օ�6N��|�8�7)��Ї:���G�jA_�p��= ؒsɳ��⡈����'ɂ_1�(2��ly[�\i�7+m||<6)i����u��y�C	�^�	8w��������<�B���Q{���2!��wn�0�e]*[:%*#����'k��GUK�Y:����w�e���
��A(����>���RAE38g���+�S/Ƿ��㯖�[�ra�ۅ2nd�>B�����1a��10����+�ڏ�֍?�R�kW;'���jW�A;�4jL���?�G6988�xS��Qdb��1���az$�^�)�]�;��lp��&v361�p���33��#�k՛�ϓ�ݡz�w�oq���!z.7",'��ɟ_X4��ঽ/�-�� n��V0�W��\S����;Z5x��>����:���hh3m��
�;"h���!y
$�j���@�:}ɠ�J�X���4cՐ���W�s�ϜR�io\7JM�h�L.뇶�$#�{�jog����p��裇|�8�$=ؐ����@Iz)s)u��`��ɍ��v��T����2kS[��^�&��a�V��7�CH#
�q T����Oo��X�7�xN�ȯ��+F�蟦�+�nmM�XݳQ�#�L!��R�_�'�:������gӨ��fW�W��}o�$n��ש�Ǚ3���f*[Ka����>�/�5f�r�̝)�����y�w�� ��Ps4�&�b�3��wY	�Ə8�ן'\��f_�Έ)�)��y��С �E>�����p�2�{{{_#cP2��I�D��?��Q|���tp QΉ�Q� m��;��"���p�Uc֜AM���c����A�s{�zn�;���
��q��q�a��Z��Er���f�:�c��l
�+cF��MMԝi�jQ_.TU�����`W��FJ}B��ঽ���w�����nG��U[7����|��E�WgG���$פ"K��me���yE�(X�P 칥��	8<^�����B��Urw)�-RX1P>nF��7�8���^b\�.6�S�Z���=��Lc�g��_oNx~��������r{�k��F�a	��nե��JP���<22�� �)�W�.�)���L6+bDi��nLϿ'��M� -���6�o�`_->P�Ou�5�,`�TL���8
#����_��mc��靬9�����z��sO�h�c|Ӵ�`<Խy�=st�%ѐ��]����6���2��V�|��B��7�� �%�g(���q��몿^9Y�M�e���Y)��[�1`	�f�W�p�s��w�K6��/�W/��n�6�[~�|�;�s��m3�=W]o��x�'r>�$""�3�C1�&0��'��d�:3�k�D�Z���K)��aA�* hy~����G����������������}�4O�#�;2��x=���Oݾ|�w�����7�\WSᔎ3�)�'�:y�e~h���jX@q��O9g���T*ɑ3hj�Dv�U!k$�o�ա�KOI��5 ���?�]V�h�鶯�S���-��42*����	[¿=)Kqu��1���MQ��[{��qXj�
�i�M_ўGw�aE�Z�����;K�un���(x�γ�>�`>~�V�)�q�Θ���;�� �o@�^�5I��\1wC�o�#�bM�g߭�4�Y����1<��R����W�_q��1W]�e������5��;-��t�W!2��� EK:��EHcNJ50Ή�r�j��·�p�������'�
��`+�}�w��r�u��,3�<�� ������/��'�A�6s2IG�(v���Q��a@��
�?��;�Q�R��W����U�P?�����I+� �
��"L!B	��A��sdj��k�Ù&�OE6��C����cf���D
��2؍�tJ��ƾy���q��B�q���,
��V�n�Gu�DRJ�@Ih����t-�>��J�M�y����A��mx#z�ݟHvYs�NsGO&|��!PE:ݼ`�^y�b��]M���uʌ(v��q���
���+h�+�+%���S��߆�yb&���:��_�4L�5��*�5��)��Q���^H�45�a7�'{�	��޸��5F�2i�(����|���B�t��W��
���+��sQ��xD�G�#�c"�Xӡ*=���W �����R���L�bql�0��-Pߙe��|c6�U��^D��AT{~s9pg�kJ@$F�*�ϯ���	�}CB��Q.c�~7N�-ȄX�.�h�h�Y_��� %�m�=m\?w��逰%fXﺌ�^:�pu���p���+���Zb<䏳�Ĩ����9�갊ݹ��1���b�wӄ������X/I���6ԛ�C�yL��-�dMv�����p|z�6��?��d���6��$vz
tM�K�]��F��0�eW8�F�Ȓ�ZU��/��z�N/����˱2ԍ녙F.�	��:~X�Y��+^�gM���U4]r<��qS��N@���*�����߱�^�b6:3-2u`m��Q>b8K'�k3W�>�.��}w�;k��}��Xδd��v�!�Q;��LpgW{�E�)���\Ť��8�i1rrr�I�k|v����r�ۻ����ϰ)1cUq`�!te�?Q�_��k�˥w����� �-����m������t��g���T�8��m�"�O����I0�
��k�L�FiY���R�9�;��=>�DC�N!��0U�H7�퇨Ža �:�2��E2w�'�e	~�lҏ]�El��C��,���x�&��s�Ro�WhTL�)cd�AŞ�{�@����]��D6�s��\�Hi�^���2kA[�������*�&{Hm�;�G��k���9����vQ��0i���r|2L�A�.� [AIROO�:���ahG�P0��8��#rLE9�����\u�W�P�ԫt�硝�7���<���h�q�>ۙ�5*`�*ָ��#K̐��3�ǔ���35^7o�e��Շ���ҶC8�Ka&E��	�"���h��U���?:Z���J���,{�O�����]I���T���/+�Q�bU���/���.�|��"�z�$�S��m�tQ]�T|��B�"kJӔױ��x�6g�����%1����S��\���Vu�:҃g�+�N�ǿ	� ���<w-���6��y����d-��M���4I`=2�h��>�+���!��ϟT]��x���oO^��U��8�⻷ ���ahY˞��VU�UA�N7�/�ՊM�N����+h�2���� ?@�u�¤P��uj&,�ŷ�yӟ�Mu9p���*�p�nH��+L�l7�yV��O��jc-�mێ~�9�Hֿ���%�;~q$޿;�m����b�s�;������F��n��wz��A�h�-���M�3v��pU��r�mj�N�ʁt�d�$���`}����#3~�V@�Ύ�R��u���|PO�9���`t�~���$��&8l�{�q7	���D�>�h�BxA�B��|��>4��+�<�?�����]M��d��t����)-��2$r

* ɞ@cd46]"+l�}�pr�_��%�L���o��+((8$���?��""Af���vS��o���rt�7��:J�N"��5�rr}:�T��X������v;�ՠ�3d���wNu�&�\�/��ԫ{S_�x�q�x�o�2�nΟ��uq�h�&�d=�(�i�C��(�AJC���������i#���[���Ư�H���]{Zv�Х7cw��to���q8��B��==Y|7=+�{��z��5x�+��pS�d��,�'z�2�o��C=����c��8O�Up2x�� ��A|$����ǂ�g��TX��	3.���g��H3{�zW/���~�oZ�7��qz�XlPd�� k�qv+�u��OR�Dd;��r��������u*��՘U���<9�1M�T�S�!�(�FmҧX��鶆�Y���=I��,%�Y+u�5�!YB��M.� �4�l�Z��\��g_���-졙�ˆ�֥M�N&�������b����䣌��L��"���?�ɱ��V�\Y�ԇ�P�<���I2����nS+�V����k�����ml׍�A@��x��E�a��F�j����~�ǌ�����.ǂʣ[� �A��j���.b(�.�3.�5��pޤ�\��'�i�oj<��,~P�Nߦ�ǫ���b��⳥6�^�ZK����F�a�p{�� ��g̈���԰a��C�2:N�"���_��YA4$�63~���g$��d���r����̦�Zt���j�%�ν��V�������t�B����@gX1p",����Q�s���1?m@����~��)Y��'��t0��I0�n漭Ĕp7u9�K���W�\Ϫ��vC�i����Τ����5P�n�U�'l �+�ö�����VOO��A�\U ��B.~a$7m���E2b�q�7��,Ch�ފ�I�i���<�"^�	NH�(���]zG�Ǎ\۟R6��H�W���6Y""<�g��k�A|0"�â��%��������6t
|
��X8L�K��x��`�K�\��ϻF}�M^��Ґ>6����=f�و"K�͸�(�ok�\A��Y�nu2ݮ�D��Y���4�=�9;Si���|B��܇S��<ʀ��n���;iᓭ���Q�]h*���,�$��;�*iʺ	�a�t�F:W�h�S�ڸ�Sp27����8��
�!kY��|2D?�,����t�������c�In�b���aX�'Ϻ��c��8L>�[����L��F��� <k��f��r��˶�T��8uT����d�dB�	" �C�>a2TW#���a��Y�#q�a3�V��r(��2��n�  rZ�:���  v!��Y<
�\��yA��@ʡn��"��1���i����0ӈ���.�,����(�Y���y�B����F'e��T������Vq��utQ�~J�]�#��yY�@	�����9I��m]�H�*��ŉ���j ?��i��Q���H/��M�!lvng�)93i��gdóJ�hy�vű�L�T�!@�1��$>��X(Ք�6���y%�Ô��w�yw~�w<r���b�=��H9���X-���M��.��.@A� �����z"�� yyޣ]��*�t���J2�8�Y3Ǘ-$�|"����>DN�@�Z˯`�ڭ`����E_Zg>|�u�-����=ͷ��:2g�=t���,�/SnA�K��b�%.�>VI���~=����Z��rh�4�0���j`6�s�u?&�?��ؽ�Ƽ�R>l?މk�Iq���z��4��P\ا�z��=E�G�Y���u����i��qsr�+���}�J���F�N�\W��f�7`� {��PJ���op^`E�+D<4�_����k�"��=d���������+>%<�E�)� 6#c�㰟D!N"��G"p]��ř;��Ε;ٌ7�*�z���1���?�-��V0��ַ�c��8D:{r-nV�q͘�E����OFĒ���ら�E��#ĩ1<������Z.,N����vvwc��^��q�'{U(u�5�A ���	-�5E2"̖(c�#e��D�-���2m�����r�N�	� �uB�0�'������DfT}��z=}�ð��(�����=s�똏ݐ��AV,�_e�?�l��p��V�,g�to��io74�>���_k�_��~���x���:o��t��5���t5wg����z�a3A��XlI�R�͈''/�R8�,	�V�3�Z��+�U'E��ϿB�#즎�R���Φ�+��-�Lה�h׍���#��z�O�.o��z�L���~iH�g3v?AWl��nIlΎA� J��%�+�ԚS�b9��vBH�!Ii�<V,K���5��z)r�~z�W�g�����7VC���R����~W��ǕB�.�Ϣ�p���1�qt�D�T�Ӏ�_#>=���j��ԙ��Y������MWVI	�U��#��d#�r��JV�IRҞ�c!^Js���`z��w�ݓ�_�rg��b9!/xѠ��C�-�.��r�Õ��Js�?O��Z�����T�:'8� ?�^�n��uc��K	ё*�Ҿ�6�ÛP�@��k@��v����
� l�͛��v� �]�_l9H���!���7���#�,�[5��()�T������UD�p ����q4n�I�@���:Z����?>0�2��2^Df�	zK�y�� �v��.Ru:e���R��߽����M>u�ǵe	��g�H�4cMs���${���%J�6jݵ�ݤ��7��������'����2^���o��Ig;�dYp�X���I�әN ���H<U���^��pL��A�K�z'%٘�3lYD��E^����H~�b�����u��7�fe��ڕ���D�qF�����I���l������9��)ԉ����h{�2O��&ӆTh����N�4���+�()tTG=�S�,�5�wq����;,��˯��Exw���n�mx������sӬ�4x)�]�OT;!���%�)`�r}
H�f����lc-���U��ܼ��Ԇ�<0����ϓ:�5/#���t�6o�
�nF�;RSr'WL����]e�֤<��B^�h'gD}�'"��L��N�ԛn�W&���~�\���|CF}�X����?�N�C��׆��d��U��A�R~/ñ5B��u�xzz��£dß������b�f�>d=5�]�Ƶr9q��_{H�Ӓ��{��D�j����w�|M`�r���L�s虨��n]G�bj��w�PAF��ǊJ���#vu�_�c�#�]g����vM|��I�+0�T��ރ���sB%u%����x�iԿ��DP�&e�w��\y��ɷ,ג��x%(�&&��.�t��2(S�<����o
�}� �� kk9 �7E֖ϗ��q�*Sc��!�L�a���9�2�.�ʏ}�;۹��S��3���g�F[y��}�A�G������`�0�lSݘ�RI��}ѩ��"��uM�jjb��U;�jQz.ꩨ�E��'�Ŕ���	/�V�C�Ez����N�#mF�);}����k��<�'�7}}��Z�8�UTTl����O���q�'*��>��?���%ì��-.��Z ����r��z��{�3AE}/���h��_
�y��&5���on��AhZJ�@$b�x ��^�Ձ���b	X6M��b�����o�]P$~2���B��C�a����Hl5~�a7�e�B>��xO�KcZd.�wDZ�k���v��$�(Z`l(�_��o-��<m-RBXC�Z?�T�w�C��G=���D�rd�R;��(=:��IbY&�M���V���H�W�=#=�����j!d| [��j>���m�N�,��}}w�c �Ӡ,p��\<�����������'����e
����@eJ��}�xFԻ{�	���ä$rƋ>Jd�̈M��������!"*J��Ptk���4v����{DN��W��Rh1Y�Yn?�5�qi��fq�ޖ�7�zz6�6	D2| �ui����L��N WU��"0����(��Ev���h����,���4c�0/?�u?�ˇ������Yʐ�ҙP0��V[��z�m���߄��K@.k���G9;�ۮ�>�m�$agR�.&�-� g}i�33�Z�N&��e���@���޽ �[�w�E�����ׇ���Oc�G,%�h�0��\7?�?�K�M*Ot�l�?��ʑ�����k��=�lpr��W�}||"�X�������W>�[����.t�����+WE	A�׉��=<x���p
vo�e����y�����l��������� +͋� ��'�f0�_(^��Ur�O!�'���%�lQ��#�~nj{k�/:��!�Sȸ�=�q�E��:g"wN|&�w�q�g(eK����C��{Tb�y��$'Τ���}�1wN�\4����(�u"�l��pC�mHB�@Ț�E�k����2��,�1@�M����`�� ��	�cy�0�c��yd�F�Ic�Z3�ؠ�kL�[0�w����E`��Q�m���W.!�����J���|n���*�$�cC΢Sm�:��Vq�U�y[�䌿"�z���b/�
x�e�T1U�!p���Ȓ��'�ΒI��������*��E�q��1��iٹ��f�y+AKK�H'!���:����r���]�B�R��ץ����}.��W��l��
�l�a��i�ɨbyQ67���i�\��q��E�"��䭭���#������NӸӧ�}�X��g<d=3\���s��B^�Aß�g b7����|��O_*O�ٰ((%f���5�V�ѦQ�sZ�]J�{~�!�XO)E�vX-"��q(��0�֬�+N�����[��v�1����6NoW���hT��N�`��!�+���nʢT�}mn,��.7��J���yޣ}�K�!t�	���a�����+2ti��?��ъO��ƌ�'�cG�Y}�ǟ��
�&᰷�S<V����
y'�6��g�{���j#�������G��xG'�Qw�5��i�w_��ӵ?�'� _Ў�畔���&6g͵��5Wyd����"l�:��:3��G!����������H!��,�~8����Z�4�)3�u��Vފ��� U�v����vQDd�� ���{*��E�%�Ћ3|�q�B\�AR�a)m!�z���R�0ų8�xm�0���F^�����z$'k�-����ץ4z�NwM{M�D���H^_�X�8�r]�	BCc�[���^�+�G�q��?b���,E �[�2������iTϵl��ͬa�ƭ.ט�[�x(~�9�
�w�N����c7�	����b��>JY_��&�|H6rv�1��#�KW�{�>�_�M*`�A����'�J���{b۶jĭ��2Vʂ���k��^y":���H�.�a����۾�or��A�'�W&��U�.q�{�� <i�G�G� pA�����7f+�LNm��BQ���J���P�"���T��K\;�V]���"Z%��4U�-j��?M��*E��5;�>4��h.0;0n���M�P|��.v��L�M)�o�w��������L��������J�^XaKTj�"�n<����[�X봸`�(�EKeOP9���\s�8~��<�����������4�o��?q�uNwe{�� q��g[�Z�=��>sΨ:�u���\�x���o���|�G� ƾ��┕m�)�Ζָ�c��.uA���vB)*�%z6p��޾����b)+b#I�lfBLo�~oc�{�D�8�P��<��Ğdn�e������r�!�~�em�7�!����ό�22���I/Ձ��`�]I֎4��:���1ɢ"N\��gj$�
��E|��H�;r�n
�]9�_�j��O�)N�OB��Q�ϻU%�����U���g�x��%b�x�d$R����1���'4ZtY�����ן��ܱ~45�	V/�)RƌM�[Z[�ٹ�O%j#�y�^ڶ��w���AO����n�\�ֻe8��Z��
�'T�iz���&H�W��QF���;��F��QT�\��]���oW�s��LĿ����v��̝U���$�7�B�+�D�O��L�Z|����wO���Ş�ٜ/�]UG�p,'�2>�^�M�omT4��lY)#���e��_��3(���f�G��;H��V���f ̪N􅁊��
o������x'�V!��?Id�����~T%Q6<���L��^�%�=V*���a߆��7;;�?�m|jp�:�^&�ζ�ެ��"��l�	�"aXe��i�h�=�o�l�N��E����m撷��$&��:g�}�a�.K���ZZ�z�^�;��ҕ�	�Żkw&����iłt�O$�\[]�t3���a s�Ǵ0���Θ0WB�[�d����U���&�n<�+ז�p�[�0�+���DR�l�I��t=|#L#� O���E/�
��-'?MBj0\��Ǵɣ�E����D�����Q�?�����}�Td�^pBdHua�R��ˢ;��_�����g*/�yT��*Z�[]�2[��aֈ�q'����(����bnR\��R���:0;<��jx��v_CW=m?V=�����"?A�%Ǻ��d�4궠^{nn�����Q���_�	������XD���"��t!�%��L�
&��<�'"(H��S zK{{%YY��GX��$pi��F��:ٛ,�t�Ϟ���ƴoq�Q�s�����)R�))����P�HK���x��i���CT�(l��*��v�e�@`-xq� (����ͪ��L�+�G�q#n����� �[F١K	UYto�W;��n
����%7�k���O2*���#�d:MBb���:��؍��~������r�;�n<��aG����U�J�׳Ԙ�:\Y�x���w�=�����[�?�^�.ʞ߈t��o�:�<2��'�}�GzK�F�X��`%r0�|T���  ϵV�R�#Ǝ���z�j�1Z�����)*�3s�t��&���o&v�G�������KO�hu|���7�P��T]�Sj��0>�M!$��������a�1�?Ѿ�RZ7� ��^eF!�y)Ƿ������5�L��u&�~�������ǃ�	̨���b�з7�H�u%eD˷���-Yt�ŀ�P�����$]�7g$��FT�ڊ�̖��c��l���N����~.��/�0�"�*�_�D�nG���AR���\ZZ��E��h���>�⦢�M�FO����2�a���ص��M�N0���_���q���+�fgm�+�[(TIho��WJ�/�L �?�<u���rG5p�	�d�U�\'��$� �l
u;�J�q�a���.���8��;�m��_Ge%T
�J/����%����0DA��B��0 �,j ��+�A�a@�#eF�ܒ��;�̩=� �FBD�����ex=*pu����$�Dp��lt^v�+??�BÝ�{1�[�R�#��EϼGDt�S��l�Y�d�0��k��VJ���Zx!��ϫ��4��Q�"P
��Msd�a����1�,�Ҿ������hQ�׵����;�d�l��N�5ip��Qsi?�?�����T$��I%������9��f���b�3y�:nC�9�;�r�
u�<��X��0i%/��k>\�뺍$F�|z��,U?�HO��-C8�nO��W��毇��g�} ��g��� ��ɥ���@�G��P$�@�T��+��S�v������h%)l�z4H�w5���N.jl9�_Tϔ[q�	\!^!��ߐD��`9J��J��-k�<q���ՕX]�S�&x���F����ީ�³�p��e�_}�#)����ʿ�D��9������n��B��8z�o� ī�$U���e+B�?�A�ɒ&���&}�Re�p�>c�3��>y��������0���7�̦�[9�^�����6��V���/��E�)ko��TF	K~i��E��J��`P�U���&쎈��k4Lx7{ޠH;��p�QA"������=��t�ǌ��sbf��f;���ǃE��v�B�4������5ho��=~��.�ij1v !�����Cl�n�����j�o �A���v���Pj]�&���Fg���(�k��&f�>�2%����� e=r	Q#�S�X��CJR��)��¿9ϳ
0?mܓJ�|W*΢&�Դ�vnix��)�r0���(b"�u�o�?����J=K[k�c�j�ޒ���9X�~k�%YU��FP#W���ݰ�������R�Y����"!!�����,><�#�E�@`nM�	�������ki�m����X�Â���+9�5��ji̢2�I���f~}���Z��M9]P�7��_�?Aj�M`��z&����c=����-���<��.%�4)��O��o��2̞*x�p������mS(����tw�o3:q�� R�'_G=�P%��Oy�pC�vio<ՍW�G�L{���G�Ö��"�M��T��c<��X�����E52�Q7�u&-w��[�����ve3W޳��3����G���yd8�^.�s��a<`��E����M*�3�1fE=�M�F��n  ��e1Sa䁶2���0J�M^�6�v�+V!_IN��U�|��n��8N1����F�}W�~�����_�z���c��>3�4����}�\��L4n�+��5t!U�#ٛ�Թ�}X�A-*`�+P�7A��}��Y�.�)�\~)��Q�̾i�˱R�!��f�-�&�U4n�,������fJJP�bW�����k��L�D��H�Y��k�3�;k%	RUsu��^��-+b���3�G�GS|�/���,`��%Š�v�:J��vO`E��J�����e �^ݦ;�pݛ!XKg=���Z�������ԕ�)2�HV���B�LG������"�����yjbG��� i�^�ڞ�:�.� lsǃ�k�\����v����iϽlW�*<s�{f�F�F-F%���T��}t[j2h��;! ϗ������G�������4����,ۧ^�,8��|�¤a#�50��;����E���VG4�_
�]��R�����ϰ�}tf�DjJ���Q7�u��p4�3S�,�p��@ ��#� ��a����m����YTX؃]�`'�VUd�q6Yc��q�7�q�a���?Q�k:�g�D�@+$�g��^pz8<��_I�P���@c�&f��I⃈ed5�ݍ�ls	;_��G󅪛�`:�� �9�E���Vހ�Y�f�歾�+�e�zTnO��f�Bu�8�8}��~}���-U�3m�vz��>�m"_~�]!݄��a�g-@` 1�B@�E���K��YbÈo�&/*��ޑ�ϭ�oKh��$zQmc�5�!���%��I4x��E���'&�q{@���;��^i<���tЬ��X2�z�7�,+�&�������H�M�A�$1}#AUK1�W�+
T�:'�s�� b�ي���#n%�5���(.�-[
����b�����)��{=�R>��
����VXIh�(޺���Y��h���-N<w��H����m�a7����?9#���R"�&]_�:��)#�e[�kb﨤���)ss��x�%g2c���V΅���_I�gΡ��QcI	�����=uA]�^����-��y�U8���Q۟��V�'O�6�>緰$0X��8��S$�~_�{@��<�C��"� �n&�p�.����m!���899���s�nV����'_���h0�ޠ�YC��C?���"+�lH�&��U��`pڝ���B[v�B[���Wլ#]D4/3̥^�/��22=y�� ��@+��~U��8wc�P��~-q\{�k{�X}J�<|�繄]�K82��ej��Sp�Q'�7Fh�����gnY�)XƷ�Mı���j����M�sW"�&����V�6.��iX[���*/�{�-��_E�5�){������6
V��D��_����M���5�_�HP���a-��_A�����������:xy�8
�1pe�G0D�����p�e����j�g%]�Ϭ.��#������̯GF�ާ#��m���,2�)RG�2Pd[%�O�x�� ��F�g������'���dc����d|��+t�P����ё���`aNN�݂�
�҄��xך�*��(�yAJ�˄3��	3?�$�H�_A_O���v��d��\1a�5��'�m���f%����T�C2e@n��d$��S���aWg9�K���G�d~TqY"z�4<Jz8}��\i�#����Ë#3��L ���J{?J����fV��\�Q����e���+7d�몦bKA�͢��)�G�{�8���exܽ�c�����ߧ���T߀0WYb5a1�.R�{��Y���e*/={��>�n��W����:9\+�UX֛�����6b���)O�9�$M�(KcI�_���Nz��ޡ�a(��%���r��E��@حIK�?v�-�k��e[����}��Ǒ��3+���ު>t��sjW�3��D���S�'��H� f�|����4"A�W�̸q���,�E��B�	��hss�����S�Ö�/�Q�y�v߭Lk���z]w���Hy�[�v�r�<����=m[�b^�b����4�ߧ��� ���6\��M�q�X���fz�l�x�p�ۑ���P0��P4d�E�n�`kf��
����G���������K2���3�L��O�;L����R�q%�|%\{e{f~��O�:�cg��h�`��	C�"���B�do�#9��?�����J:�r���2f����~�ʧ�;|�݆�k]-�A��O�Vĝ���t���w�m��)�$�E|ϕ,��J��5�_��)�L����gP���v���l�.�z!/���h�k��w�	�P$�o6M��"W_WYXvK�t0_稐ix��ȔAUyT$�=�V^l0�ֵ��u� ��wΠzn�EpP�w�!�*�K����s�=5���a�n�I�:G��%�/c�,�ܾnI���(`���{h������f{&{"������1�0�/����D��	�=���]@��� 4�&H7ߟ�^x�N�-��+hnz'g�R��n�P+}���	�o�ѧ���O��u�����a�bo��5RQ7+KQ�_���x+M�La"�i�������?���vD����e�bh���d
?���@���ڭք�ߛ��0�8��,P��W\��wTH5�g~�/�)Zz����3C�o�-��1a`�ҧ��x?��O�	;ZO�=JG��<wP��9��4��gP��J��R/�1����{��e�+�^�N�{�'��O�e����0�-���{�(+չ	?}x������Y*��+��z�e�9P�t�RN5Q��k(��⬟�������v.F�h��ň`�a���� ��U� xT^�����*�����`
aR�,�n�h^8�H7����/}����(����4ī�%���W�d��1w�-Ƞ.ɵ5�z�7�}.1[\�gM���W��ˤ�����;y�Cֲn4V�~_5[�+�HIo� �b�K&����kr��-C��xա��U&m2�FF�bE�J_��c��2�|!֣E�*O�8����u��a�3\.����((,T�-[J������(���8I]�q���DUJ��������d���扆J������f���u5�)����}U�Z��V��чt���L�d��6�s�"�V���'�<���v��YDp�oEѿrP�o��ˈ����K\�.�ʒ\e�HO���e:�JF�>�l�tX���Eg\���K��)���r���hK�`�W�^-���� ��������z|�(lRZ�)��,}�	Y����gĹ�+#���!~s���ᓠ���6��K5޳��ffo�j=z�E���p"�b键�s�ŕ����$����g2!�e��_���1!�>��>_�%�+.,,<�wП�B�������>>�1��+{6�hۧÌ�p�?u�|Ѝ�Ho�ꍸ�H\w@�ȧ�	�6>K��|^�j�������[!o��Dqh᲎����t���v2�~F�{xs�v��k��%p�:PW��
!m/.`_oXS�a�~	� ^�Xߚ��gϋ7���Ԅ������x��۾y��Zk�S4�0c��8P=���Z2��]S��H s45�X�V����H\+̥&�'����!^A�R��0�r��cU
ITE2�����&u*�-v�F�y*��*2`?�L�Y� 7��V|CS!<IUk5��68�F%4L��lG�۷���'	����6��O���:��<x�u���g܏]6���=/���,��"�:C��	߱��Lڋ�lNu�"�?�d���`7�L�M��j���,���@�{�<��3��'|edaR��[0g�W��c z�a�H��VI�8yu4?���j���q��#���ց�
��su1���o�&)�v�������>Sc���O=��>�f��٣E*�uI@���G
D���,Am5�4B���L*�?���d��h����}���VZ��[�%G�c]�i�U/ѯ}���6�/ >�e�0���9Ҡ${�W�1#x���TǪV�@�5��GU������e���}ϖ�ዓ�9$]:7�-d�#��;uc�=>��u��]C�jV�[N�<�ԝ �P�H����϶SKK,0�7by�k�yhO�[�,�gh��BQ�ѽ��Qt9�u8F��7Z����)�SPsO����mk+�S<�;��E�������iQǘߌ�o(R�o�g,ԍp ��M���H k�������kK"�ZnC�4�Dw��Q�l�B���K��F�R�3�\������,*`�׵Y��+1\�4����D�3�΀��2M�Y!^����ͣ�=֠��l���Fz�l�ݳ\V��ս�����`.�i���<��1�T=�'��dk��bظ���r'�X��3�gfDT�m���-S_�x����ǜ�t� ~�6����2�m�P�ʕ��}����������  ��瀇�	�����[�E�=�ò.JH#-��]
��% �K�(�tIwww+��H
(�y/~?�����G<���3q]3sf�,`���U��L!V�S�U�^lv�SE�&Zf��ط�nc�`�� s��H�WLYbӒ;�}̊5�s��S�4 ���Cf
��Y�T����ϭj�A]��-J��P�cQ��C^�li|�
��Ra1����#r�^������֭*�ww.e���ʛ�TԾ.2m)"L_�6ӤhM�Ԝr�.Q�����7KRhn��4�j{�{	'U;`mX�p:�����5eZB�73����(E��F	����BBB���,�7�;[[!��<��ld��8O|_r��R;+&��F����(n�l;�tJ接x��~x��(c`��ʽ9�ׄ��&
6F�e��Й�9�dӶ���೧Um7Թ�����cu$��H�e-�懢����gժh����Z�Ko���S�l��$����E��(��F��$�ly)����/�9�ڒ��@�~>V�j!HR�;������.�CA8O)4��l�L�0��wne��2999�����d-�@1?:ӥ����]���o�w���5����%�fk����3Α���ƹ�<��G��!.�gO�%�_� �=
�ɝ�v��v��p�4�3`6^�9���M�m#�3`ʴf��n�#�IK�4>�r7Xj��N�'��J�睹��	XX)t����XM�04�ܪT@���3_r����5p6ו)�X��� �ĺ����E�v�C|Q[@]'��)��&r���1kl��d��s6U��8�U�A�BL��H��[n�qͅ
�ůe�x��s���V����7�%H���u6_ϥo��޼�0v�d�mD��]r�Q��'9S�l�*a�^����Y��'8��������P�&{�>� BrX+j[��2�HA]|_;7�bѣ�0c�df,��9/}3%�zXP �TT�$�����Sk9�4��t�v{'�F���U�����3$�%��\����kh9zˊ1C����67#��g)bȽ� �U=%�X�e��\�����������˪>��N\G_XOWf�X�z	fK�Nd�����KZ�o��>$���iͻ�� }ڡ�?�\6���Q+�˙N��Kۈ� Ʒ��߁��������9��p�bE�ǻ9=+V�nF�W��BC�VH&̪;�f��g���=y�ư^�����N��1f;�k���:I&�i2ӹ�_��h�d8��e"E���	d�X�^�J���G@.�F�b1,_I�io���̝��S��ڑ��%,����_���Unx,� �d�U�����1Dɶ���~�Z�k����'4�e���Cqb"8ưѵO��c�5�T	�ڝB��Z��s>�`�G%�6
̬��f[�-�S��,S�D��&���0�������H��Z����葃:5�����	��޻Q'�u2�{�ۣ-��R$@k 3�!�,�Q&h��
��A�%�	��:��@f����l�04�r�߅�ޘ��܍����þ�&��n���#���%s��徺��d<��m��˾�[}��ꃆ}��w�lJ��
��w��*~��߃f
�H�ҳ�Rbm�Z'�ꄟ��bVs��d��fE�k#3��{r3
�]*U�t���,�	���i�^��88����#��^�ܭ�#Y����,R��]c��"�=���eL�K< ��-���G��?n���4(�����0JaLN�̄�G�GL��^��I?����c�����M�9�N��Y:h�:h8���>�{����!cgx�'X���_ZMݚT�'�ܐxk�`K�l�!3΂��-�36l����]��Cǌ���a�T�nj���^��Վ��w|5�����	6��P�ո����i���W~^5�yw8w䰳�Ij��М�4�G�L�PGfg�?68`dr�MXP��t���'�|�R�%��=�=�d䕌dKpL�%����?�3DD3�����;e�M Q��q�	[�IkY����>�#��ƭC?�b'Kg�y�p]������l��᾽����U��t�D��c�aO��2�į������tɵ�ϔ�b;ux9�?h�Lm�L��+UZrV���������U���E�g�)��'_�0�]��P��Z�����9[����\�PdR�������B�t����,�a�Q�FQNP�궇��>��HᾸ(�4���@��sY��O�mK����J���`t|g!1��{&�p(Êq�o��`�t���_������m��� 1DM$�\�P�~�#�{2�X�T�ac���=]{�&c��8)��h�+����"�z�����^%�Z<�c�"i�����b���o�-X�����=/������qc�Rzq����܁������F�Q�3�
�r����=���̠uNV�>�4�)q�����?�Y1�`��u`������8ӸZ�~���/J�׺�ߢ���ĝ�����Y'�)E��z-Z��k��
��t�a�N�k��bN��	����Mh�����7~��w-~�-P9r@^�2�9���A�=^�N�{j�5L���E�R1H8Z?�����xm���zl�����A�+�g3�m,�E	�^�=�b�fae������*�8a�(ʳ�d?��:t���l1��C�� IE�{�y"L<N��8z�2�N�/�l��göO�N��B|�(��>�0]�%]l|z߹;#�wІ�ڕ��o�-�li�\GD@�V����0�@��l��u��N���6q������ڹŀy�Rܱ˗F�B�B���(��h̍	J������Oڋ����y�sR�;��O��9ƫ(2���OT1W����_��B~�`f�/�9ԃ�����Km#n��R�9f@���=	&������EL�Av�<9��D&� �|i���.�{5D�����Ta�o�LY���oįA�r���aB27}��`[O��nm�~��<N��j&���DTNeg��Ք���qт M�UW��L��*��ã��R!�A�$�����f3��=��A,Y�̳gO|?ﵶn$�=x.D��%��R���ᣧX�ܱ[�M�[�v\�zh�P�	���E ��{�fK�'-5ō���#�\���
��_{m�~���ں<p�+��ì<Ǉ����^��r%�n�d�|�p��j�|�U��\�$�[b�����t9�\�
���Ĉ`�G׺��z;}.´p
�{
m���CꩠZ~� ��C��Cf�9��CBB@0��YYs,��G�� 6$��)T�{*��%iI�ʭd���K�LG��
�U���t0�Y�Ɍ�t4]�;�q�*�׀p]ꩻW����1�.�_�S��&��0~�� ���O4`ŮpK��*X�������ʲg`�Q����1��Ϥr�$��|�Z�=���=�M��A�@+e�ED��1��q�� �)_�X{d�E%##H�q?%��ĹA>��F�V��MF�ԡ���l;�-��T2��QO�2���X���Ϭc�U���Ώ�&��2ܻ<�]C,�02fD���o��bs�w��^7v�=��D	NJ�*vt���]N�}���m����	 �ɸ�G�4�]��p۴�3u�&(����V8��k�$N�%����^�X��]}���JW���.�s�#`}%U����p�mS(�w�����
�����S'V�ՎZZ�4s��}�/d�>�I�2?�!�&���E����z�m#���#�!XI��ؔ���qO�}��I5Bۯy$��7���){�~D���i6�k.�K]TO3�4����j!��T��E� �2�=ĶeM�;9S�Js�?�L<RFNN���羦�{1R�������~h7..nX�Jޛ{/���  �"�����&`)4���ܺl��"!���t҄�Wu�]�;�������҅���'D��> ��ѵQIK�J����~�ۊ�3�P��甪���gπ��T��m��y0V�D�"�i�!�eˤ�!�u����Ф<JH���tF�Q����QS�ϟ�-~BP�R���d2���Ng�eW��l�6	(sZ
mkJ&\U�l�Pϵ��9c��f���u���
��3�3@��Z&��k�y�)��|=@�͚�����Ǘ�kym��N'�LPYP0~I�7@fc��I�һ�N΄6�|)�α���_:�B.�?�����(�9���t��X/Ʒ^�� qBġ}>���q��p~ڽ�P�o׬A�!�Цw_$��lM.*Nʛ�'�N4�n�ty�i�%��IHHB;)�` k>�����I�,$���6>�'	T��l��|�����Z ���׷"�6��u��.��PN �65;;�� �l�=��D�&,�{vg���D1Q��9�X9�'hB�gwZ�
��Wc��vH<�V�9��*��y�f	A�s�.�#����*�S�jIEK�cY�v(�YQN���?�9^1�sx.��������>37w�)�mU���F���S�GK�6	`��N3���նi����!�O�餉e�ݠ�x�H��k>f���X��b#Tj�� ����J��0�;%W]1K��)]���}a���O��{�sSe�����րR=N��q�L�}{�D�Ç |���3�ݿ��܇���F�����*Ձ)�� Z����^KF����n`+Zw@;#����R)�(���+�	�^��6�j�!�0�w�r��@��H��k��Q��sJs[��ϲ��Ƽպ�B��@� c�6�Л�x�g��ܟ��)���&��p�{
���E�t>Q��&^I�57���3pHf�J@l�/ѿ����}�*� �P���ABƃ@|�v094���+V�&A���+�q)��"#o��R��L^�n����i�;�v�|0,�,"Hq���(��v�\�<)���7���L#g}�ȝ�#]�����1	<-���w�8(�9Ce����jao�xm��8�lzm��ǒ��B��eB|��N���Lf�V&7�`���a{7�`��$錫oi�{�i��}i,���1�W�p�t�粁_}��^@��ˏ|+h��t����<���_��V0r���(A��>��$�B�cybe�e�����I�ZG��)�"�Y)��K]۩9Q��O�՜�~�!���q��Յ�� �zV G�U1STxH��,���u�<�aS	54gSvR�G�"4+�Q[���X�P璬Gy�����Ҩ���efx�+ӑ&@%�F����2�)���n2�1m��^�"�ބ���`�z�Tm�*��U@�X�d�Q�^Q���Ԯ��{C
�?�z��^BfW%(��k�w'�;�:�O�U�$�߸y�Y�!�w1�`5T�-���t�A���2�&p%"��ٗ�t�&�C�4�oj60U
�[*#�]7`jQOOkH���O��j#�δY���46O��-��hkF�5���6H��p�۳7��R1��'��O炨Q��R�91J#M�IF`z���~�K,�7�%��x��)��\�`�Qr�_W��(���kԘ�#�͛75�^�tia�C�c�7a��KFI��� j���C�@('�����(p��%��o�g֭��&�mP�]{O��P7�y{qpp�i��O�?�'�g��1ܜ,qI�5�섛�,���X���!�Jd�9�@���O~7r����i�U���l{�ø����Z��襛]�d��|����t�_�W�<u�!�I)5;�]!ݝ��%u;!v�4²��^�(������|��`��W#�Ll)�8��^_Q#&�_O�x����]1j�#\�J��<ߍ�,|��~��r�=�7��e6���r�K�WY�W��Ѫ84��!�a���O֯���#�3���U���Q7Mm��	 �����1���j >�o��K������ʭ���.=����݈�%�Vt P���^��r��V�_X��vJ[�-g�z'�^Y�W�6��5��<ק׽�>"6-��,e�@�b�C���t��C�,B�XAG@�*��I�0�i1=�)�f���s�ý6���q�������IV;�z;H��f��j��s�~K� UZx�κ�1*iw�*�D�K��.F�t|0�����C&�����/z*mTҮ��4�ܖN�#ח��C4�2�֥���L���E�Q!H��a�)Sh �ˡVz�T�=�<2�	�����J�~7"���T��k����<���s:��^�!6J�n�(��As��⮕z���*<�z�.h ��L��_�-O0�͈ª�XE�Ӓ�jDٕ�P*J�����h�|Wh��h@�g�<���;+N����4���4����G�Q4iB�7�ɛ1V�a���h�p�t\����h�H:Z�p5fu���%���~��D\�J��QɆ\��7�%<>X�_<���l'G�w�Qq	O������_�� tAly�]W����O����~�Ģ��|����qp)y`ً�u]���3'�.����eq}Oxo'ۂ�������H	���S�Q/�l	u�v�NT)m��)���҃6��x�����biG�z]�8F�{�������Y���`[��HV����ێ���67��Yw�n�$�鴾��C�i�r�}�7Djn>'�&��Vy
�}��>��'����5���+,�(H�#�F�/��R0u�����q�"��΄�R%���v.�W1\��E�-�f�A�,<4 *ȚTgF}��<@R��P�̖u�0\N�f,��wި��ֳ��3���c[U����fVV*b�Ջn�+͢�QF2��nI����jw�� �$����}4�*y�K���7E���f�"�A���Qn0�$�Z�k�1�#���^NG��rU�F�_5x��V ���4���?<���}�3�/He9<��T���ỳl�b�u�3D�|��7/Y0����^��)������[�'�Yk�C�uuGk�\��ܶB,�߉0��``s�Ka��)�b���Ƀ��PP��Q|����zb�u���v�U�P�T���[���h 5X�p���4t�c7qy���
�T�:}��?���LOR������fkN�����k��Z��E6��!�\�Y(�Sb�f~M�<�'�o��t},������ǻCz���ǔ�t{�c�+�/j�m�*�À�-D��+�>Z��c%�{�j}��r!����l�ި�8��D���;�:aA�y�?���7��A2y�/%�;0b`�X&9E�=f
0��`wHY�Y�S���������'��MOQ�}c���h$�佉+)��ۨ������L���:�yc�d�˜$\*j�S���q����HW��{�����{���So��Kt�.ƅ���"a"�%.;NH���ny��E�l�c�O��R�=*W��
��1�>*�;a�E�@��w)��7����4�ѿC,���f�j!R�.��ݓ̹�[c���v�Hɩm$ex�ʛ_�¦	�{(=v��27��r�I��.�VQ؇g^��� a����~��uT:��ѹRj\^���
Q��6�����nQ��C�n�Ol[����ƚ~�VT��ҿ���
��ŝ;�-�3�kvu��;2���e,hm�fK�"(�-��^��ӄq�9�ǿx�% B���+E���N���1�}~����.��Tg�yL@i�la�m������������z��g��7/�Q�K���V�m�h$:>ܑg�8�6�<h�U����\�������Gޤ�F=����t&�$E�S�3�义ɲ���>�!��DK8��!�����l�{��qc�3
 �����x��nA4���Ǭ�f@%�����u��V���`��Z��XZ*?~l$W��6;7G!	��-U|��A�P������xL}8ABg��-nW$ NQA����A���/ֻ����� 6i�J���j ��F�?�jң���xm��j3������L
��noи�Ͽ��Ѥ� �q�/KQ�Q���6���8G���^C�>B�]��>Ńd`�IIIQ���=[�u�@��($#�=�`��I�L.]�75�X��G�����R1�	��2��K��y[5Z������6�h��W��f�E���~��d�~����ݽb�7��34�cB<¹��Ij+�3�V��͘T�K���e�'�}_��o{�6؝�yx�������Xb������󼹫�<���������&&��,^��ڇ�m�1����]�K�\C�����6��r韧�KR�V=�j�a����FBd�����!��׎���ZY��(D<HHH0�>!��qf�wp�k��F��e,9_�-a�E,���o�2=��*9�p+ɼ�����	Vp|R�ꯈw& �ߍW#��ot�1O;�n��K�����е�}����}lg�I��������!ψ��(=�2�]��Ơ���ni[n,�zU���q�ґ�t�l�c��"!?���-�j�P�gJ�9�A��)	m���������.�YMƚ.w�K��f��dۂ)�}Z�ٷ���;t'*�I�H�+��Dcm������俦�_O`3��H�,��!~u��c�k�2� �K�[�8Zt}/�Ec���ݡ?錓Chϰ�k��^��_�o%�����z���cWI����x����|}j�W_Q��HL
F��&z��Ɔl�E�&�-#&������ ��} ��{�] ��k��,m08ߒB� T�Y9�|�c�vd�uL�[��_eb��|�x%��:��z#_�i~~������X��m�rI������[��_~	Ƃ����\��)�k����ro�]U�)ŗkWQ��\u�������^�<�K�ϵ�����}�E�>}�� ~v$r���mdo0Y_�&�N�_�0���4�ŘH���SpBQ ����N�A�,0����r}��~UL�����/ZBi�6�9O(sJdJ�����C(�2�/L?��}v�<�����\�ku������糙O����	A|'��o�,e0>(tǮ�$�Zk���Q�_	j�|b�i��پH�</J����A(P���J_f�MW�f+��Oǔc;�����'���͑��z���k;[����!�tkG)/:�x��ČA��#��)�C�1��n��f3��_xET�G��b����K�c;n9��ފ��0ml��궁��O���hI���'�7�t͗��W��|��i�NI���D�DG�{��,�߄���LEu ��"y�w�"*��#Ux�
�^�03�����u�.��􉌣���Dz�^gb���V���ۻl���㏐�	�\X�����cv��������'xc�]f�]Bmɀ�6jо/��e'�)%B�VR���tg �x@�tc>�+��sT�<J��+N������D,$44A#�|�T��}�{s�ﺵ�I5�3�_��*A�XE��"y�%>>��-d���3��2=9��{����ۣ�\��'���umM]��Z�t)k���YvSt�oT�M���V�[{�,�b�K�m�f�0��Nhh�^�tz��l��M��~�Z^<S����={\�a�>m(�����w���prrbM_�`����oF��V���607c�!��{w����]?=u����<d��P�җב�"���v����}R���4�`c&J.`�WW+��};Kq9�x.��+�Eu��j6A]�vf������] �S\r�w�V��һ���Wa��>�@��Lm�C��]���F&���2�T�cl������s\V�����0dt,����Di6`gU�._6���\���Dp�M-ɩ���i��B744lu��nL\&i�B��IhvRB
��(G���47h\\S�JL߻�R��1��2_5���%��J`mzS�sK:3������ >�m�4���$��(t|�7��&��\��ac�؋n�v6�?�@y�A��'�tbNT����/y����bk��3�x[$��DȽ����a��x�_<�)_N��L� >��n���bџb�lY�,�/�����Z~p�����m]�;�F�]�}��D��fVb�'�8�]s��B꥓��땛�\{!�x=�Y�w!4�ch%�������N<���i�^�C���^����cIc#�נ��L�
�m;�P�\�8����GT\\L��F���v�ύ�\�W����\!D>�]O�:�`��~	��ϋ�3]���j����YD�K�������"����^��oE5�I0І���gU-�&��Dnv��M�7�X�2�ʳ�
5��U�%a�������rD���z3�^�����'&.��;��F���v��7wK;�&�����r�p����pjQ�-Ś 2��f1ck^չ�ݮԩ�p������a�r-or*$L~b��"������(eRh�g�`�C�p��.����o_���lh�#3� ���m�W>iî=t*a��A�
�ӁO�ɕQǺN�����En�I��bqR��O(�⧾��)�I��α����@��,��]��8vyT�w@�X�'H�!�2�w&'^B���F>��#|!
[�݅XW�bM�������v��cgO`IU��i���*,��w�Jg+@,0:g�T`,�#~8u�>�E��=�ѭS������Q���]r5�]�G����և	"���OUX���!��nz�4�`��Ru���	�J��ͬ��Je���h,K�xo��-~)�q̷H����KP�_�}���|��݀8����1=���+ۋX�D�f�vȧrj���*�>���&v��:4i���$m�W6� ^z�d�S�J�WD���B�5�-]���и5�e�k��\e%��e$L����}G�~;Y���R��ﴷh)
����/þY�P��T�rkޏ2Lg:D��.(�n��N�kBP_�w�ĒV��1"»����M��_�٩�����!Ƌ��
m������%�����������e��I�r�M���z��Y�qZ��}�������1�M0�m�]m�g�P��XS�g��}D��,�"H�:\#o9h��
$cvwwO�������D=�xa�����߃���};;��kR,�n����S/&`�=��~��"3nn|���hn`�m$�-��`�<a҂��|u�m�_4��p�y���=���gh���c�ϵ=��/�)m��b��B�6^Z\���]b��4ˆ[`����?������E�{} /5�(�dh�Z^0C]��J��6-�30�
C�����aX�w��y���`���$ۏ������+8Ecs�0iKAd)4n��y��Ҳ�@�#�����݅��B�'E��UI.Uы���wZ*�n�ak�Tj��J�V�'������&��4�7{ܐ2ZCο,%=��5��-��Ԯ%���V��g1�!�� F�� v�yl��FQ��q9JR~NX��Xo�]52q!����c��'6N�@o�{�.�k����w�530� uz��ї����K|�����Qٛ��4�#��^���}.N���at�4�ޜۓU�+�v||��E�i!������#*YD&�C��O4Z"�y�c�����,e�3���O�����d4g��p:��݆{�p;�Co��^~r���9�۞Ω��b���m_C��Ȏ'���>�.���Ѝ��I���������V"E=P����@+��Ũђ�L�0��`����KE&dbQ�2ƿ�g�3=H�vЎ6A��]�꭛�p�b�=��w��Lv9{M���Z$���o�������*���hn"G������%~�\���ӵ! �Ȏ>�8����M��| ��~#g؇���f[�YN]>$��!�M4r���.W|�z���f��^���3������d��o��m;[��l�Z�9������	�ttJ!t�:[��ۭ�blpuL[�4o����ɕ���L<#C���ۄї���s�<]���,+-!�			J�Ǔ�8�EZh�Z�,&LZPC�c�1�ɇG�34p4�;Y�畗�(Q��Ur���-^]�@�&,��*������jKY*���M\�8���;i9uvgr�1,k}����ԃU$�|�ڸ�9y���3�tȔ���������I��:��ɭ��n~�#c�@��_��fmM(���k�h�:�Y�Oo�?Hš��H�`�������6��0t�J��t?��{x����k�8J���7d��V���:;F��W�b�����ެH����XZ��ų��T.��FC2�!�nv���6 PE��)ۗkN�-�
w�u��H�4�0QB@@H)�mEY�+�[�ow��*(b�`��?�&B���.q��� ׻����QM`+�@�X�a-�V��d���Z�u|��[�P�5���mД�=�?���*�6W��\H�����~�5����@�_r.���p��FҢ��)<���lzX'	���57�ji��wi,�J�q��4���������]�ʽ?���?�:u�F1Vx�v�VY�.b�oL�շ�i�';l)!nQ���4�^o�"{b1�|�?���m���)@/��|��g��I5̗�W��G�&t�e�? Icf5�B�S#,��<��/�^4c�P��;� Wd��O�K�9璘�M:*Ǝ���o����H^x�Mp�)f,:>�'�G�ނ3�FF �Bt��9j���M�w����<bт�d��c�J
�^��|@�@�����:u{�dӎ���.�j�	�6�׌�֣E�}�}��n�\�;n0�ι3�i��e+آ'C�GҺi��XȒf!�G1�r�Q3��M��}
$���R��ȳ,J%Ô�&i�!�R!z9L�Bo<��B?Ԇ-r�,���d0�̃O�9<�
��	<\C���C'�����"�~V��Aztf���п�찤�tHou��(7��l=�A�|λ�XU[[X�i��.E�1tH/�[x,�1��������������Y�ڗS,�g��߷�Re8"#X 0�bi�E��o�fGS��4��W_�D�Q&�f|��e���i�2��Q��#���l�ᡉ�Yf^p��^=/E\
wYk�i�+����������侸sET7�>��J��,�v .B��G]-N�[=�;���ďf����OB[${�]������V���8у����� �3�輿�[{��cq��O�x��`F^��ۛ ���?RpId�F����)��ӄ/f�e�R�0�>�18ȹs����,�����
���¶@������_�����3)~���G����W4w�3�V3	�?�sܓ7�S�t�o�Z��~�!�_-�m�N��cW�nǑ��ܜ�O�Ժo�SO�� ���і�<����_Q!;@��6!=���ͣ=����#����^����U��L0��Q��Iܑ�\EHQے��� �sM�w(3�-��L.%^/p��'�%��A H%D��y��B�8�G�u�u3V�dj��V���S�9r�
�`a!��Y�n	_;Pz�v%��٪���*F��xR��MgX�i^����`|(��j� �Z�y�K=�� ���n�٘K��ć��e�a.�0F�\��6���蕋��)\uXP���"9Wz�.vu�U66,�	���>�.��|/������L�����6�����Ek'���kډ���%�#�C�:�j�LQ��zF��R{��eV�,)�i�x��'���"L�Bw3�6C&��t�ϒ��A\��"��;���v�غ`,�;��.k�]�H#Kge�뚥�<lo��d��>�;��ϛ���_�G�0�'l����=�q4{s�ب�<I�g��'�&��v�Gr�QAf�0�MGǾ뭱��q�m�w���>��^<) �[}>��
���u�YV�1uDt��#�z��Z���u�L�3�]�!Ru.�U�-�˹Gn�����SNj�ᠽ3,��G��Ȩ"c���^�8�0��.��z��Ơ�6r��!�B�c_�S{�qQz�'�}�N��9���cj&�X��-��i�L������-f��L�� �n[���Z~O7�Ʋ� �v���Un������������g��.'�V$�����5��K�q�	.UM�i��л?<uX��'V��\^�y��Bg%�Ã���<���0*oŔ�`��-O�o��\������~�5Ao�a�^�j��
>K�����K��	{��갨���ӹ����Hn����?��V5%0��#<Zl	��Ή��V��~6r�3��Sf��[�)m�M�8�����������kߩ�9��e׷����+�QB���
þ�]��@V!�7�$����Ha��9�B4��k�ۢU<<<~�W�P9vv�IC?��j�u�F͔��� ����T��v5	�&{d�U	
��fѻy��^	EC����%���*�SJ�,�S����s	p��;�!tΥ���A���=�O���"�]�7;��O.�����f��N ���|$����!�8gg��%L��Z��w=��=�uZ�0�b��pg�mF*�R.[W�8j�}Ey戵���v=�k��q��p�8j%��Їo!>���� ��V��eb��:����u�HQ����
-�iP�v^��^��+����0c���h!�D#��M|����OA3_��9��n�].�$r�FO��x��{��d'T��_9W�l�k�0g��ϵL)�sXu������B6O�� �p�EB�54�³E{6��GRb%�{0��M��w�W��7�%�	¨��Ò1�f^PpU�0��K��o���:e�n�?ݳH)r�̸^%���.�Z?~�5ۀ� JW~ܩG��T�|�xrr��Zvm��	V̏��� �'��&��:�^��O�3�Fi��z��1�U�d����ݏ����o��Yr�	x����N�h��@�ow�L�Y���xG�o���+�oڷ�p�!����)+YM�لZ�>#1��~0��=̽�:^�^��@Ƒ�L5��t�~��n�[dV�G��c �)|>�����'\��;�Et� �=�{��0�ݻ�`��]��'z�V�.'����Zi.}eS����H5�+�ɕ�:��� ���i�(����t����g	�����3(Y��x�&mUhS�CGdނ#��N�O�7߫b�Eo���UνB4��x�:�ÿ[ߗ� �_X@o�݉0�ie�q��� �%S��GtQrpZ	>1pn���_#���[�+�1�7���wu+̧�2�ߪv���f��x,�IB�>����X�K�l��$Y��
2�3�"�z�ڄ�2�&H.��('��W�4��%lp��h����t�V�������̓�{�,�b~~�Ɍ�֪����~̀��yS
>�L"�r��)�}�B3��bC���/����qm�>�o��d�wᮽ�t�u_���#�3���{4~�����G�%m��)Z���D��.�1�s5J�c��]jg�L�����H'Ӛz����(��&�����lL���A!�F7��I�Gzzp^��KN��^Ճ�b����S�b9��l���&-�NWs�x'c:����Q���v ����\4��S&�1�su��]�.]�/�C�j����Ą�@k����@�c����#�+';���9>y��¶�ٜ��jPoÙ5:Kz���gڕ���c��{f4����C��LU��MM]��LE�O{▛Z��v�տ���Ψ��L��@�K�'4S!����h��W���:��VRG0��k�b�<%����O�Wkjj
��6*!g��7/�f�lJ�7N�񎼌O妹�K2&�0���*������"y�d�����J5Z`'�,F�--�~�"���_���� ݑ�ʍ���b��Gw�&����W?g��G�+]sg|o������2Y��Faݜ�V;g�t�0�D���<��hg:�S-1Y<�Y��c��$������ݲ�����ɣ�d�n���g6�7g��I��~Y��:O8�GPs���ǥ{��a`�擊q-X98��vJ�HCa��.�y�1�5��b#O�匙>��AL�m#�ֈ��8�8΍�s2c�����S��J �a�n��Հ��q��cC�n�4:ꞟZ��Qݼ���ڹ�e��3�"��q���g����e��x7F����-�7��*�ޙmVn/�M�MvЏ�7Jvu[�p���>äiP10�Um�ژ�4	�n=:����P��Z`/�D����_ ,p��r�q��l���W�10�gg��2d�z�|!��3�as�E��d�����r|||]��V&zM���ۿ)Q��ey.��������g�[)�X���sU�o=.)����cJ~���m���L-&����B��Ń�H��v�M\���<�_1�7|[��ɵ�=
'!���!��(o��ރ���X��o2
��Ռ�S��r�\N:^�Μ���/)��%a�� �|*�<z����#Y"�YZ���J� ���^�;�F���>Oΰ�mgH�4ML:�d�?���d��Ì��-kS�J�t�Ċ(p윝�|�	�Srk��>a�n�4��X��S����qdV<D)6(V+��C�3]���^���+dJ��J��ޅҷ_���ג2m�V�b�[�%0���1c=Η�igAf+b	���N��?�-��J�<�;F#�k�N�Z������5�	�ق��6y�~3�JXp�z�ݑ}�L��d�y�a���H��=��E���ۋ.*�����~G��)+-����~{�7���G����=y��E,&�VX�6<���[h�)Y�nts��m5k�"�h_ؽJ�������51��	w2F��{$�G���t�[���zэ:����qK���i�:��/J�j1�ªƓ9��K�g)tp�{�<.����y�T���H�'x���1z�=�	1���^����V�oJ/Q�����F��rU���ɚS�ݿ�t�t�S��(gl\l�+H������su_����m�m�c��j2��+�=�YM�^��������g/t��Y�Yپ�}{�U)t�<mngٟ�	*?�$����kb����,}䨠q۷"4zd��4~��g��yzT�b�
�%,՟e��C�l麋��h�W30h������g�jB� ^]ڏ,�5��kc@+�f���S�"������cMZ�ىv�&�ޤ������[ۖq����CZB���iiDD�AJ��A��S��:�O<��?���{���/�.�����Ŏ�د�/ɞ���h�D����ǹM��?v>��F0��Q�pAt�5��s+�c�� �_p�G�,�5L���p�P�*Grn�Y�;S��E�q��|��bI|@�c���2o�]��g,�MF��=u�ae���0-(�L�����^A��̹�����T�'tT��j�)����wciY�H)<A�&�3�� �Y$;Isp��)�ؾ���fۭ��W�c[[[�F%-����_Zz���B}o�Ů"w�����M{3^���	]�Ѯws���n1'�
��t&��Bv��*������c��}�\=�6��,�9�{,Lsϓ*�g���-��{)|�D��|1M'�S�pA��N��$$�	�l�^g,����]�E�ڸ���%�4��gO�oT���+����w3W�s�A�G"UN)��t|S�"���õe��
#?L�'0���u�[[������IHHpv7�#\�C_��Є'���G��q�r������,�sC��3tց0�7{����3��"]����,���%2�'A��X��������	��A���;��f/��Wލ�cR�nA�B�j�t�V9RU��d8� @u���;{2�7���7A�'��*��@'�#��T:�8����G�iq$.6ؿHC`Ⱥ�p��Zپ�K�Z�0ޞd(��4��A�/L�D4��R�9r�jBLHP����0˙��uPؖ��vן�e�=4�ϣ��.K�M���}h�a�W�[��6����U����Պ�N��#8�)�G�����Gz�D��a\���jii��1�cO�1R�E�_�� ���|~�������T)#�K���x���=9<T�r=���_)O�僷�	�����	#��6+�q�L�"@HT���Sh�Z��$N��;w�#]]�n���t�Ⴖ����ʡ�F���C�	���7-Cx<{7��m.���|ŭ|O><�Oy�r�)oY�Q>o#N�4��+A˾�j}?HbЙ��>����9�_���=f��5bE��3���O�����te�����_6�\X-��NNN�oK:���Չ��,��s*�"�
Њ��0Z	q�#g�
��"(}������$"��2�ں:¨�)�c�HT�!%�+l�ř��jLV�		��;(���=v$)�e��#��x��������@Z������+Ŵ����҇LE����~㟌Agm����4�%$�i¹]�����ņ�>��~1��ڠ(�O�9�.$f�V^o�i1<K������3�}M��IU^/�Wof+v�t�F�TMG­�7��-�P�"�QO��앋��Α�a���/Y4I"���h��P�)w�n�u������d�l)�V[�#qUzh�e����f�� �|����ȜW�1��z4�_;��c��E.��	G��.)b����6�,��( dg23B�6�w�A�O�&�r�)�W]�A�Dr;)G)|����~T@< ���x��-ʁ��R�`[�6�D������vA��Kղ��e�hs/D�	n�.nh|�l��A��L��\��Xf�軞(t���&�S��n��jH�;.YMg�vرo]�ni27�/��i�
ߞ�T���3���)k�y0��)�����}��������B;�w�'h���6J>~�&�I���������`WD�Lx�,�V�;�D���sRR�tK&\�q0\n��S.|N��/s"���R<�1���W19)������t�߾&!�%��̬i��U(r��(�y:�M9m�6v��v���h���
n(�50��),��r��]@�/����8��z�g��4���J��zg�/�7���P��(�W)�P��J~�8w6��xFD��3ì����ڠT!^�GI�˸��['a�4�mo�J%!nQ'm���yo��Z��_/9� �t��N�%M�%	*9�V~�p�>ɟ�`�	7����4
p|ټ|�xgK��3�ʹ����W���a���!��m}}=�r{^�X��-�����R.��ke�`j��z�l�'="������u�z�_~JG��i�W���<�f��pC���.��%�[�^t����A��l�?-��������J������nư�ȑtط�������n�������?���>(Fo��ܨ�f�+l��ݍ��Γ�)	�ٶ-D�ow�6|O����W��w����;�6<'�YT�q�/Y)��i0�	�ݘ���tb���WE��'ߦ/����;y����6Iľz���#i�Wp��08��8�U\,��^���+��.���K��>"�w4���%e8}���{d��X�a7���`�{NG���0�h]��h�Z` >	|yW���e��U���q7c`&Y�Ǐ{>=�����*e(�߿�x�_�����������}-y��]BY_�-5�!,���U(\+��meF��ťV�X���<��ddn�%�M9.���O�5��'�Z:B�0�~	i����b*�E^�)��o�H��CJ�k�3�_�Yi�c@8%�1�Y�g����b�e��M|I�1C��l�К��=oɁ┇���>��eB����*���'D�y>ʀSix��y�
��'Z��ѼN#'�W��u��eQ�Aԅ�G+��ʷ�o�;-^��	jB��~I����Qk�TTX�Y��h�d�����9�g��3Y4񬬑�&x��;�;$R:~��"<�����~ٴ��gI�:+F����d�lkml<����>��i����^��q�8r��m�h�g+e�Yąa��(9��C��$M�n���TY�.�qi.@��6���Z2�ٹzl���W@����-������ࠦ i)�W 6��_U�st�[)n�n��su h�O��w�
���+�*�Y�<ěE(�/�\K�2@Q%��D%�����~��eQ1�$r�G�M6٠��M[[�x���\��e[��UH�Ae#���u3���� aP��Ǒ��i�{}��3���ق��P���P��O�C΂�Yh��K���j� T\����S<&�g�g@jEӮ����^�P�crYH�-`cҷ�ˆm��l]r���D�9�^�*CL&Q�s����b�����$Z7r��^^��ݥ�cc�������P��BՖ�����o��o�����ʑ'
5������,E!�����Xn<7
�|��eJ�ۄ'5���\@Q�na�Fb!ҳ�
Nk���K-�E�r6�N���T�n��/
\���O�ؘyJ/֎'�����!���~xx(�6�0?��o=ȵw:��G��w�p�ŀܰ����K��	������++�3�~�3�fvRJ�ţ���D�H���Hp��%/��)��9�D�}�E:�ā���M����fe���I�&bO�:�?0ax4��A6F�%���[��v�u.�)AС�����Q�MÉb|ċ��n�����Lm`?@
h��^�^Mf8�3�B��LFrQ`)|���<��`�ɝ��iT�|wkKI�j}�vZ�Q��P���4I���������)�j�����G�T$oE�ZG$�6��ʻ�iPꊌⵉ��X�$��@8���n�D9	K-ɸե��;����)TTn�C�*��@��q��*mm�8{��`q�j����S�2=ݗ��x} �/Jሯ���r��o5[�W}��ms{� �T���t����c�At1�uD��(PiTB	{ܖ�xA�����[�5���j��L���x�w^�6��4�pN��Kl�,�v2��>����r
�[�p�m�(�Y��g�X���7�gEi��9J�4��E�"��.��6�1nq�	I/
7T|���s	�^�Ъϱ�>�ܕ�GX R�4���p@o�����F���*�f�#��5,mT.}�)�*��g�\��p`�>�D���˫����{F
�� �Ǵ�U¹�:�$��ٍP�������:�y��ŵD��YHQWmBe#j޾In�H�|8��ðZ�+*��C�#ѻ���j~��۠��ǣ�U[_��Tk�م�
�T��kL�p�Y���M.���,y�k�,�D�n��<0 ��C{i*����G0�i��I�Xx���3��P������?������אq6�[�K*�x�sjxJX��"� ����<�O8l�H�<�ؿ���23��q����|NM�w
ц/��_���:E���P��@T���af�b��b����U.T}��JM	�J�p5�.T���~�ө<��H����4�' �m���k��k�M�}_��OÇ��:�oF���I}i�`���� ׃��N���4`���!6',}����]]�|�<V~���3` �Xݍ�ꂶi~�����tS�ˣ�	�ѳ��wM�F:>��o�"��$Sv+��͟f��&
�5�o���'*_ǲ��К��/�y�����O��4�)TF$_�񭱊���¸�����I�P�#Έu����_�GͪK��T��A<��.�p���\WS۾<��H�`CKF��Vg�>Q�y?�c�T��ķ?��tmW:�6�(8;���;�mxG��)z�����ㇱN>۾�B���m�B�㼘���Q��N��6ڐn�w�N�f�ۭ�l=5s�8�T��޷��͍���f�4G�]�~�A^�:���88|U�X��K���' 鯛4m�����f��5y,�^���՞��������V���Q�����������<�+�	��^l_����<f�L����s��HD`�Xl���.NNSW��F�����K.�]l-����Lx��
)��[C�Cr���>Ɍ��yC�蛝}�dDV��x�|��N��=Pa�l#��V�2=���Ϗ�^�C<�,��u̕�瑗����_��Ēr�R�?U��[Üihi�#/���4u��;���\?���bb��ɲ�}���t��k��}������'��{3FlN�s/��_��K�:�'�}�y�#^I�e��R㍝��#�Y4.�E	��]n%HN��t�=�L���!Z�d��Ί� X�Fl��W�K����6��8���R@ \�X��K<�����nPD�@�z��H�Y��ڥ-�{���t�E���ߌ�g�<!Y���r�E�&���@ iCp�'�eyGy%����E���7��E��� ������~��0�^��PD��Z��%j�{X�.⤈��v�T�8����=��ĳus�<�����^�P���!�Q;���<;2\����1���ž&��dH�Z϶l������7���ȟ�}��o�˘8T�|���$"z{]�0�7R댉=��E���[ϳ��}����b�P�S:����T���N*��+9xg�۶�V�x�k=97�w,Ufp*Õ�J���;�3��\x4:`�G��P�?��Iڠ�M&nW�z�v���1�hkl��_b؋�~��*M㎨	�W/��S����«~���m���b8���~\Q���G�K
����9�1ڔ�%z�Wg��W~X��`����V��{���hmJI�����A��]O�R��o�-���B=���`��(��CM�<�@f��ej�������^�0^��0���.V�Z���u�c+�$7R�p���w��V��եQ�<�츁P]or���׿Z)�R�{o��Y���t�oI)��-����3S�S�WD6�0�~ݢ���������Luy����T��3��G@�9@��#��~Ijћٵ�AI�(����.�-����Ǐ��7"�����o�[�x����'s���:�������XkeHSh9M��}�y�:���ȪZv��W�u���w�6#mӃ�m����l(�CߵvΔS���Yi�GՏ"�c3��^(W_ή쫡��HL^��\I$����aĄ��@����wę����v���<"��Aɍ$���qPoI�ڧf��ͫ�=<<��o�~&�鯑��$-�U��w�%\]�o���&�3������F~���~
�A����u�����U�s��x��}���#@��(6HU���Wz��W��bKf�@��5�>\,�l�vO�ψ���qTh���vw"���5��	6�7�/c����q���L�ߥ�$����1>�ԫk|n�KU���"��9�}���拥v�'��aǁ�ȿ	���Q�0B�>VAL��(�1�?�c��l�`�(De�ܣ���7oG���X'h?}3���S�զK/�$��	tWrف%��A"���'.=�2ŹF��4�u��(Q=�^�q��Y��=Ԅ]���YY�x�L��S��1}yY��#ĦJ���:��Ҫ�g�/�6�r�k��"�*{-�?p�wS�p%!kZ4����%%�?ږ&���DA��c~S'����P� }���r�D�N�Ƽu*Ґ+-�������^�b�<�Sa��\����"��E�(�F,$3O4xIHs�9��ʦ'�e㧅�t��q}���c�J���?υ+U���0_Ɵ?Ǣ����Z9���+��6�Lz�	R��� �9��� �n7��.�U|��|�Mԥ[�N�����a�_*X��x�L��Vo��n�d����ҞxN���] ߆��.��;Qj�E���������#�G���=�垈�}D�bP��҉�=�t�rB�Ɩ�rDx<t77E�o&�m�5
=��3 ��/d .��BN�����������s/8t���ܗ�	:�����7�n�Z�l|�|����x.��~cc*�7�G��t�e����Iǹ�R�U, �) ���$�����cߘ����Da��V�L���ؠ+O]��N]x��AJUY/	�.�U�闼J��`��&�x`��g�L���t׆���2,o�`)f1�t&Mh�{{��9x1Y�8��i����+�J��	�M4��GR<����Cg	M��e�.S�}ֳ!e��8>>���X����v��w�1��gS�:H��BR���qQA���#,��U�|�*�᩹an�jl3��R9YW�e\��(�������e�Ĺ�D��D������|ё�3N.�<����W8��!4��8�j�@被O���0n���l5-���r vu/j�$M�@$&?�G���y����fJ��(#����v��t�ŏb����=���L�QD
�l�12M��|���Zr��|���>��3�'�Ҩq�2��<�p@ܳ�)ډ� �~t�_���P �Y�����(VD����n䠳��`q�R{���e�n�Jkbr.��2}���(w�@ ("��V�hh�zq� ����z<�y�Z���(�3@�����8j(�n%7����,�IXa�r�/p��`{���B��,�'����\�ʳ{�� �u �P� ���^�^x畱�R�=��Vj�Mju+[�:N,���!��!^�!4ש��GO�nX��9�%�b��ͫ�0!��m�'�b�TS�Y�k5.�6�m<�a-�,�k�D 5�/�H�4JZZ%~8�׉pܿ�J�6ZC�Ё.�U#�����'��Oڶ��z��a��z?��Y
��$N X'��¯�#��)�U(�7Ӓ�;��3
�3M�AԺ�� ���P�	�p[����n�r��*��&F>��:���	��F"M�h����\N!�����"����)�8_D�&�~k�h�t�L/��	1n߂��js�R�ς\k�e8�8�Hd
Z��_��u=V
��Ąs@�m�_떻M�j\�lTt�"hR��ۼ`�V����kl2<�SY�_:�����v�F����KX�o�%�+�ϛ�{?��;XU�\��ö	l��b�&YQ�%'J��TM��)+�w��G�*C��<5�"{L*+\D���~�-�s�֒ߖ.=Sʨ��Qd�(Z4�L"L^zA�K�ԅyQ�����6�?���2p���r��g'4���2Ew�<���±�(��y�h�VW�����'�):\���?�湯%^��O�iŲ��
�dEǷu����m�PL���C1�/�����t�6>�9�N���難G�5���@(6�����yYT,Mc�=;7Wt��J��O��$;T�rI0U=?u�v����{��k�n俕�/��?�:OL��@�p��H�,ҙ[Gɦ�]״�������=}�-9�!���w��5
�\=�\��>^�o1��6����/
�__��R�">�T��RU��yb�qMcZ�~WuӼ�m�i�8.�қyJ��qt��%;�;L{�эFCiڦP�MN�q�y�����mK�,쭭�>!W��bg��B�!]_n��ػ�q+�.Ur(Ce����sGmcR�����O��ќ����.Ι��{㞏��}�e�V��C����㗯zP.s�9v��xX��(���\���[�-����N@� ��)'K�P����m��r��އة��m���n���\����KH�BH�:zgE��_:p�������D�K�A���+�L�ѕ\�:����#����@<�"�G�(Ж�'�X���ī�덱~�g:qp�,%-����wt�ms�^�,�d8G	�Dg�V7ߧ0�qԐ�ܔ�Q��ل�8>ߒIN��)�SUU�6�.��*�������e�H�����XO��$���HP ��!m���mJ�Zc!7P;3 ٻ��F%�pS��~������� �ɤƾ`צVS���O%�P�!�-t��M�8ҖW��R�U��I�dJ^c�M�V�n*���k"O�C�����l"`�}]Bc����\�'T�ꬍ���`#�'{���y��U3�����^���?%��E�l壖bI�ƿ��\��	�H�:���ӿ]�0�#������F�����储��y�`'ح�f���u����
3�
 ��Vna��Ǉ��į
2pb�x��XS�V��m�$*����k�a)J6�U��=�ӂ�^/^�*ZJ4G��8j�;��[�*%ԇ0�~��c�0�~���y�<���]|�:i۫zX[_O����_�-���*�Q)<���uϕ���z�\��*[��mZ�!(�a<�n��NG�K�v��d��I���a!O"Z�{�� �]t�"s�S*]��\�͂��G�'+Xܨ]9�m}b�E���L�8��0I��ի�sy2n`�[���d�R,�O{ۿ�,
P�0���<��I�4OX�fN$E��MH���lK�Ol����+�kaQަlT]D��B�)����� ��3g���Y^�����F��8����</ܞ�W�Ws�R|���_=sO�J�$�9��ໂ�!���q���X#w���3��QT��zҘuj�l�A-^u�wRu\�����e���R��ޫM��M�-�M������3�^�p�<	M�߼���Z�V�0��� >����%J��?}I�m��9+L���3�s�A:��!�,V�����-�a��8����u�1�Z&����w�xVUwo�w��e��@d�r��=�nV�k�\���ɩ���7�M�yi�>�6�.C�>�U���渨)�bT *���}�����ːhR2��nI@	X���l�lm��)T=�sS�o;9y;@�)�������=y�AJz�Y�K9w_P�׽咸+uB�� xxx��{��޶�k���5�h�'�Ny!^�Q���!��.Ka���N�����>~O��l��(��ϯ#!Y�L�c���Of�Ԕmll�f}��e-hq0�z���**�|��:��owI+�h]R�HH���}���{8}yZ���JO���}�:S7T�^k-��f��HK��֢j�v�V�� �`q�j>ĥHjuiiإBX�!���N��V���u\Y&�B��
w�o{��z ��0H���(�g�r�w�ծ_��u��<'W17?�s���-'�<<266;%��y�#H�+�ۼ+��u怎���`Wv���I�](�
d粝k$�a�~ �Ԋ[�o�n3��CHo/w���vڬ���ϴ�A`i��G�����F�� 	�'HZ�WڗQ���?=Ȟb`�f�eb�Q=�U�s�q&bj �����*TqCgu�Me+�>���
[�i����`��'Ml���ɨ�U#w�����\�q�.�j�>�ڡ�Y�7���R�$��\�>�b'P��))��ev���%N$��Q�
�.}�_B��y�6��䌝B�J�j��v��/+9�E�Vma��;���)�xm��>0�<Z��3W��3�����K���AEX�Eg֘�b�9⻩�����y/��M�}�볲(ʛPL�fm�k��=�ӏ�=[G<����f$0
�V�e< ���[y�	ҵ�� D �]P��P }	�ߚ�ٽUR�(�X�kc�\�F��a�?�20x�q1�ͯ�LS�jf���8��19��/{n�g�da��vi�<\)����c����te���o�3k{=�V��鳬�ݙ_�I��*oOOOO9u��|gl;�6�}5E����=��|�'X�.g=ex�y� ���C4Y �����*����QX,wf�g3��^��q�����
0�h1�d\���:
�m����.YD��V9�U��/�Z�®H�f��B���St!.9]��!���$���]��?e|MO��MsZ�i�,1����X�;�Q��eʞ\��3�0'̦mD'ШL�m��2���G��-5w�̩W{C������y>t`|=n�:Jc����,#�X^>!j�[�~F����� ��%��tq+R��	�N�m7eLk�oǬ����K{?E��v>&���4b$�f�2$N-�)��ɵ>�� ⟙�(Kjw���+��w�������uU�����1ǖ���$�EGIU��aǂ����0F�B������x��GWQ�{ �[�7A��eg���T�1�Җx;�{���
OT~���)��0ǫ������ch�-D�?[G���o��ӉaMY�� ;:ęy�Z~Y)��u댿�
��8nF�K�rvd%�E]�fͬ�XL�*B.p��!��p_|�o�re�0Ȣɴv�C'ٌ9�b(!aJË�jgeBf �#)�8Jl'�򩩩����;�=�TtAi���V��0�Z�L���ŝ���Mdqd�ko
y��?�����N��Ts)2���,V?�?� ��u�>���P�C�v�Adu8B	�r�b���3-y�����*|#�Z�s� �D S��ue���2]�]�4�\]B�5<��!��א���(�Ly&�ز��LE.�����cQC8^́��t���q�c�1guMk�^d��5	��xQ]�uK+��w�����ƈu{�@�X���lʭ���5LDv:T����cޖ ���^����]'�i�c2��� 5H� �urҨ���;s��]��]����eQ�E$��S�F��N�E������%m�>&�p�B���Or	��gg�C�(+� �e�9����m�x����QҢ�`����b�Ω3�C�I�?���k����]_����T�;�ҏ5�ԥ���y���K�X������׌�{�Ɨ����&d"d	����Z�ꋃ�eOo��B�X�)Y7�[���l��+����@Y�@����$�m|��?I���T���O�$��(U�<q�u�j�/-��$Ҭ�)�R�z#ZЬR0)޻C��%<z�#�}O�#���c���4�8�n�y��&�j�n� Z����^�ƿ���,Y�L�+�(���N���&p4C�Ԇ�a���&��L�صd���w�F�r��Avd7Զ���,�L�o9@;������4�2�����y�4�Ԛ�%}l�OÛ�v9,Ӭ��r�3c�����O���Z&�@��P�Dx��I�E���G�~H��+����kwɻ	aa)�8@w����~/N^�tp��njx��6n�
rA�>���L���v����Am�b�_�æu�r���Q�h��3N��A@��m�9}�<s7���㵳���={���Bh�y9�_i�d�����*瓏p����5�/-^SAY_,L���D]ˠ?�l�����N]	R�W=P���t�g�������[>�1�o8�\z�E����'ކ��53��!%[A�n�*�9��}��;u�iD��^Rfxn#T�Y���#�^c+�Zq��1[K#��y���fim� G��,A욆I��>Sva���]r��o*?,�d�Ǎ;�9���X"�ơv���U/�����D�C]���f~"��ӆmg;D���[ޫ5ﻗ���Z4����j�k4�}{5������r�����v�|��آe�t�{�\��3P�|@˹��Uʎ�FY���"*\�g���RQ]�L�!B����'�y�UNn΋�݅;o�@Ѯ���6��J�@Yb��QD���	uu�$$�f���a�9��W�^��)ޮ�	�A4~�>]r�uPz�?���4�0[~�E�uzg�f�E������m�揽���z�1���V25@�H�6�T�厂;"n����=
H�O�W>�l���w	4N���-r��p��wz8Ih�8�އ5�a�|��٫�bv��M*��-�c�i�*�S����	D��!����N+���`�/�$@�1�U_�L9+���q�kg�'��6�������m^��TJ(��Al��8��|K�O%��L*`���Z�ˣ�x|���c6���Ӱ��o�e趤�~����� �������V����x,��NN��w�� ?
FM�[���1�����P����)#rH�O@���)�J�cخTlm�:*��F���z�G^X�W<_�z�]v;ċgY"iL�O�j�>�������p���qw���\�w�{�X���ȝ&H=���lJ�j��T�x��i�L4�QZ�\^_�C>��f$Tn�u];k�_���}*���RM�/��s^�O}`ތ9�^J&�8��{�:S6,�㑨�\�@]R)�B�s���l�ϳ_���zn�o�������Ev8C@g𾭧F0�����JsUF�9Vw�O}9M$#|ww�"�T;uJĩ���O1N�
C<u*��Wѧ��FJG'5���u������M*3����8��|J9R� ��R���h�M=�����::��U!%��o�`�
`x0���x]:2�
;�<Ps��o���[T�[��r�9]7�k/%�sj[�Z=���/m�
�v�"�Y����0z¯c[t�
��^o�L
Uw*@�ؗ�N޻�:�@(]�1f��뮵z�P1e��?���q �06>�j���B����;N/-��]�7��[Q�	���N����/���KYF"���k��=9�l�$�K��@lj/?��m��$`��)��о�<�b8v��f��v1}
�['����c�R�G��X�P�N\�t��������J?\� ��p��Z��1t�:���#��ީ����fu���� ���0783��C��i3o#����nC�ӂU���o\�t�Q�ߗ%�#�&a��vc|�[N��FQ����w�:��x��ׇR�#0�^�P�l��DʨN� u�f�y�!�x�+�WX��e��)�DTڅ�����on�6��.|ե�"�B��S�cDr]z�c������4��r���
co	>���H�+E�Z/��������Ȫ���**T_H��#��y�T�]h\өH�q0`ĩ2�εi�����T�6�xp�i��J$�?`������'b�{A§>sHU��R{�iӛ���j)�f�޳����s�oy;�Nz�q�M6�Ki�36�4�6ʮzŋ[Y/�����i�����g>.�p�@G�劖�]�*@�ɇ�G�9�b��02x�:������a�I;�rN��ɘ[�>��3�HXJ��N�t��k;}���͐��$�S(v�~>?���k:cN,��3���h�"���hbWC�:�y���7߾3�M�7�T��=]�>O��;�O�5W }��%g((E⺭[�U�
������o����^(+��tG�;�����~����B���O`x�4u��%7W|c0yU΢���'od�[oԨ%�1�ʱ��b�o��1������O�'r߲ؤ�k�=Pf��p#�.x�6�4^��Dķ*n�0�!���E*�~-��ޛˎ?rA?���k&�9�HNv�?�BGr�٦,6�'Q� <-қ�B(#!L���~�m�"^)�ޣ��j�"��T�;����J�̆�����4s��D�ƈӉ��q*׺L����e�_ ����HNќ��y/�&N2�j�6��Q���E��4xΧU��3�w�$�	~���Y����K����{L]���4�|���Qb�.��[�`��6a6\�dﾫ�~��y�����i���.��j
��8>6k�g���KX�F���9T��&8�8�����{{{�ȫ���5%��g��� ��rs�.҈[yb�^.�L0�ܤQㆅL�L�̎{�B�|��_�S�c�ȭ�*Vu~��-��6
;v�4j��ˁ����`��}�����/��O
FCgo[��H��_��g��3y���y��&Sp�Auc����ψt�>p�9""����:�]�8Kz���`�r���s�ӎLLP�����0	�nI�t�سmm��g���U#K˂�o�u������W�>ڼb�95+�H�h�����̕��߃�>Ɍ�2ݶU���jP�v|ƾ�&����l���"���&�!��u���Џo�{�8���<��ޚ�Z������iUm��%"�0DZc8J��%z{L��A)�%X�u��c��G>�(c,�#�t����wMh#��H���]g~����3{*�s�@�oedkk�)�J�+��ч篼vʄ:�t�,r***�p����R�L�;�X�z�kL�q��X�d��x��6�" cP.JH��<����፝*�b�.2_�k��
�M�7�Q���-��26��b�+���|8�o�:%�xw%Ƴ�Mq[w!d�`On8�Rf �ч����f3�����"�/`C-ʦ�ԭ��շ�CӬ��ꧮ��獘7u��xzNFQ���b�p�la��x�6�ͦ6�.'�����{�i�Us㍵G`�r�I����Q?o�w��AȘ`�����㦵�(���Y���w�A���5`@Njpz�3�� 	dc�1�^'U$	l����%��F�ޤ_yl�K�w�6]�V���{�'��ּOn]�(`f���϶��i�0|:�p�+U����&�ѽ� �W4m�J9�1BU{B�#�7��F��a8��cO�=%���l�q�c��0!� �>���*��XD�T]�4��N�zK�����ڣu�І�Iz�������\�~�q�h�wX�&����ss�_��7�_��Жš��	�$��z��{���d�������"ls�H	���Ȗs���@AF��cI�'ᘮ��B�Ѭ�xj�Em��>Bךoe��0
*�˰o\�����I��1�������M���a�=uE��",��r��E��A���˄?*���E�D>�?�>c݊�s\@ix`�5�G��K��5]7�B�`��δ��v�t-5�!^W�b�#�]�4�&ح7���N�eW�2K����(���8�@�<Yp��; 9�lXHO�@Mǀz&���j=�t�a��[��5��b��C�$U�svfC�XbOB^���<��4�y4Kd������}�p�//L��7��?��4�����ʾQ<����{i�z�P�3�t��L��c����)��_�`9�#?�[t��%�)��) ���/{2����I�i ���P�v`g��O��X|"%�'�g<X�g(l��J��6︬�Z���?��E�,���ð�*��'��fK'���+��s����C���%���N��h�]�r\�[i�t�+�R߸�+ ���9��;n\!���X�6�"�@�~�us��&ŢqlDs�p�Kj����m;Ϲ��o���Or�0|+:��I[��!��vt�<8�@��UB�T�G	A�A+`�^� ���,L|bbU"U��	�-́���/o��DVR�+�r��l��$]*�\�~�̗�ݖ���ܰ�#hhud��F��Oko�l���y�tߏ�2�BXS��o���J��z �qf^6��m{��$e��d�
���5�=�%{����x�~�2��U��g-3q~P�<�\ay�u��vf0y��oNj�e��fTV��>����+,���=Md�#	�E�z�@���B���$�Az�����'�#��p��&r�M��߱��k�������nʗvRRN�C��D��&K1d.�@���r)���,��f�*��࡞#݉l���@�oO��v~�����l��S/]�@����j F����u��z�u��\�b`��)*4z�o&�"��?"�"ֈ>%D�n�pp;�	l���-}��_fr���&E�EP4,�d��}V��xz�����Y����.���C���]-2+��\�a�ծ�m�ej= z�)���@���@�fb�R3�dmwW�6U�u�T_�
U�����KK,ͬ��ZY$��K�rQ��m�ڱ�5U6d1�U�������1�*�P;�`�K���r�]�0l�����!1�L��>�s��.b���K\[���`_�N�~T���#"����!��r�g��z�?��6��TT��3�gޔ �p�w��_A��$?������L�5��S�f��؇|	
N�}�^�5����]���ӆ�q�L������P;��1i��n��~U_B�~���'�Ly���ӭ�����}�����l�\C�'�7]��
���/EX�S��E��|sPF��]���?Ŋ�$8$#t"�)[ۺ�_�`i���{�\]����`P�7©('n���.�ck:�6"�Y=*��<�pRą%+��ҟ�c�_���榁��C7+E�QfH�+��{��L�C�Q��;�ȍ!Sv��+)Q
���)��P��$h�%3��-�_;�����G %��X���6%}�S������C�\H����%$sӶm:�S��|9 ���kʍ���(�:��L��)�[�8�X׍M'�d��z�Zʶ�ۤ��f�%��}�K�-�-�?ItKd�������k�:�}����3^��']�a�-^�qf���鯪�ϝ�._.�%;�t������9]��_�mj�\�w��}uXT_׶���� !-�"!ҥ�! �� ݡJ�t*��-�1tÀt004|g|���^����ǹfgf�Y{�{�k��q\������ �T���܌���z���/����{�+�O���/|%�\[�-�|���T�	p�>�A������*��f����;(a�n{���,*�#]� KN��ˤc�,�'�yg ��)ѱwM����xXLz�G��u�ꝕ3E����3N�)5���������q��˗3��n� >�Ƚ&.�\t{�	�_�%��{h�r���n˹�m�:}� �}�࠳@�F�c1�ss!�};B���9s��u���C���d+A%����Y\�6Qf5����JK�>hß����ق%���?K�氁�d���viA�@F=��I��az�qTgpC%N������Nǋ�cyq\�q8�ZS�ϴ^?L�MM��Ծ�=(��NU;97K�JXI��w�I�J������*s�49��S���-I�)��NC� D��CI���0A��T�Ь��H����g6��{���t�}�ٴ�*�^����8��c��\2�z
���U�۟i���2�Y5���8ǐ��������0�O�8��L�`�yUn1�u[`�஫�ͦ5�󓃽O	���if19yL)X@crr��o�}�ҫ?�h�1A��M9p����i��%G'��@ Pa1g�qK�`c�Ɓ{ǰ����]�=���z�dC"C�y�������U���1�o����f��E����N�d�W,H��)��>� ��ټ����>��������єV�/��&�'W<9If[!�pEo��RBP�{.��P�x>z��K�7���[=�ho]-�5��gX�`E��?� ){nj�N���EG
Д2����'�5�pJ�˽L�|'P�h��F���8w͛������l��
V�%LLV�j޸?G!��V+1���S_ ��7��7�����5��r��W�e�#�oދ�.�3�ȭ�&QN{�{`3CCk���4�T4CkS������^,�?�_���\M��[qxG��3e���w�|�$��Z�@Ժ�5gS�tK�5���Kآ`���b�3Ȣ�wѤ�"���@,vܮxL{r�d���I�kй��0�S
`��"�~��˕�~&�X!_U:�NS�k��|I��6���^�.m�nS��CF;_n4�����e�
2i�To��Bj@nݜ(mj�9�,�X*M=��q����T��f9Y&�X#��]�&��ŵ�Tr���/���y'%���M�-MF��=�Τ!����Md	�i[' 1h��g���x��������P�S�D���h<�[Txz_�^'���z^��.]x9	Ao�k�hc��P^n|�HMr��a �ٻ�D����6�Gv4�Y��o���"
��d��|�v(�)�T�j4o�iL�j_�Z�m�� e�2	������;�V�M���N����/U�����?���Tea�r���h�]'Mla��3++Ǌ7�I�M�n��� 4�[RM�8�äTTbݴ*��G�e?R�|K��|��Y!��W:mo��������fq|�_����e(t�I$e�����8�mcA� x
~7���Jo�������.�
f�T��	F
����.Ȭ���@:��>$״�G>@�H;u~��+����NFW\/�Dɋ�ܗ]��.�}G���j�Ѹ�C�˙�ۃ��^��k6�kF{�,Q��~�n�'���I���7u�m��I��ؿ������2uщC*�z�1�}OE�*�l�.k:���Ζ���Ҕ��`y$+�K���gffo����*��[���?�%\��{��.���E^�4������n�rzi��p��
N�S0H���1���¿�eۛ�ֻ�M6��{&�Nߖ�l��Yq;�+��_VtD�s��qi�3hi��lR�^�'bi�vm-�o��>�^�c�����%^\��t�"y��C))���ɲ��'	K��:�#r�����&S�f��ں�n/�ڤ3��ۯ����ď�n/J@�~ߦ=���x	��j�{BP�dk�u��J_��)��Ykཽ������J^��;��7��(�N�mn�Rr2-Oۃ�U�2�M��)�:���>�@΃*\6���+�r�i[��	>Ǥ��,��<����H1ԁ$**BJ�`�C����:o��ű059x�����M��*c�ø��ht�I�zSR�:+�(C�,�z`�äl����Lz{�}У�3������G��.S�"_��S�}ЖNnl-�xXý����]�3�3��+_�����4�M�a�n�[�Y���7~oDg@K�/�֐�l��Y�{0D#�0�n�7*�i�zn��%'P}!l�<E2#R��`���eu5�W1Y�%�u��� 5r��=('A	�dL�c����vf��7I�g���}����S��k�3�6����Pȯ����]���5�՛S��.�Q-��R��z+j1�RXlR�+a�����-��e���
^c�/��D�n�M���6A������{�L$V���@w�C!1z�ˆؠEZ��e��
�'j�}�PYA	m�)�uH�W�`Sb�{��[���{��:ld���6�|�DE�h���Vd؂4x��x8���(�~�\��3�m�o�_�n���.���������	�Q�1da�R��?Ү s��� �#��At��Z�	��100п�759��'�l`�t�c��q_̳z���QF��B��˩�_�Sp�j�3�+���p��Λ�^�9F���|��Y�	��o		�U짡��Jn�W�;����A��锤x�v�f�����Q�s���-��_�<+`Ǯ��&�Kׇ:�$��u{�޲+K�X�\��r�Ș#�rZ úg��<>�*RoQ͇�<?aY�p�;j5N�|��`�/ܓ��+g�K��LnNP�$��W�u��{#t��M�f��0��V���u���j1����66�&��>�$��7��>Q�$���L��.���WlʼMV����(B'�\MN�ϯ*)�BL�oqٙ%Xt!��^a��%Ի�{cz=�i'5�8�8��OS�L���S�꾹��_�?�xr��V���Q�v�	fh$W���<"��ԠJ�0[��!���%'��;Q�^g��I�3���ͮ5#z�Ւ'h�{�0�����F
�.�3����yHyV;�O�حsa�#���6��j����ig��y�[�����ZYb���{p�4������������V&fOx���Vև4��J9�d�LTj�W����8x�T?P5z�����W�A˖G<�������g�=�t�9?t���+�/����x�3�yE2�O#
|�6v@[ҀSd��{�8p��J�_���o[�a�F�u��;wS�K\����N���!,RV�:���B,H�=d>J�h���b�� �Eq=�tہ��\������h��q|xl/���93K�)���*���ͧ�.�.n�GKM�������1� ��O�!�
Ty*�1���γc���sS��RW�k�&�����r���<�2mR�K�o�/��E��ƽ����yG�����.���l�)n��T�� v�I�0�r����/��N'�q�0�
��[IS���4]苬�},��@�:�L.�ڃI/�O��R��zPqyI�/AJ�܇'cݺo��
�n��qP#Y�RBc�7���U7��_��� ��Ϯ^���m���4م>���(��y�gX�N�wÆ���:���!���)�c{B�xb;����e����,���̭�"*�H$���������FV��B�45��~�<��;��q�0��~��͍l�����K�౟���R�s^�d�=Z�B�O.<�Ι�q��:N�ʓ�k�nO�9$˛3(Rf,_��0�ݹ	��Ԥ����E����[/BQr>�Z�i�L'��|����{��x�6Pi|v�����z�s/p�~���V���������լ��(�5�>n����3���@r�ˈ�?#��F�W���a�f�깘�OZ\�W�bOoj�\GX�ט������|U���I��x5�4K�dt��	BuRl��h�lw"V�0�7�Z�Wt'lbM���s��!�t3D)��5uqyV�t����|�����~���p�x����ގ�O��������d� n���S `��ABW�����L�_H̃5����fK&�M�X�������]����7�\_�uTi?�$���yU��H�뉸~����N�u3+��-�i�X�Zn{Q6�[l�]�������ۼ��N��r���Ȯ��Ղت��uѹ�f���P����0=��3�8+6�}�z����󮕵u�z�o
|�>�"��C�`SA�>v_6�J0��J'����G�]ƶ�ͥ�^*��O�NE�v��2�h����٧�C7��^����ݞ�V���H���F٬�~6��Rf�^����9��6m!��nm�R*Ă�<�ϗi55�o[O����Ӊ?)$~�q7������sX9c۶��}-{rpCے)�4 d"��P�c�u���F�&�6�f���������s�v�ܬ^�В"HG�z�L�����7��g֩6��z��;Pln֘Ю��gW���+����d���r<��v��E��d1�,c�yӵE:���I��O���v�h�&��Dx��1��z�!��x6v�B���yO�Icf�&8݄*���X{���U�������@f��$�֔�С�)"*)�gK�b$��|��g�D�#;�'�����(A�,G�q�m�^Ǟ�R��t��suc�K�$��#������N�0w�<����e�0�g1�m^P)X��vZ+O���k|z	}�7�r�_SJjG�=\�F�C��{�W�V!��-Z�"Ts�Î�^��v�)���t��(������r��,�f)��;�\�H�`�Č��Y�	b���M'm���GiS��ب��B�>x$$/��� ͙�u�\���J��a2�f:|8�*T��W4OX��{�J�j\�?��U��|��ZƄ&����I"�_�Db�-��2�\������N�W�
��I�Ĺ�ܠ#�m��D�_Z��.f9�3�4�������>Az��g�&(ѿY�<!Q�)ܚ`�t�l}s���<�r
[����[][�e�765�h���I�	/:��w,%���R����^���)�!9o8��h1�@�_��}r���drke
�o��g�����S��)��{8c�S�B�h;}8�6^�38�]������i�/X� }e1��;\7@�r�#c:XE��~��lN��ŤN��ʷ�5}R���YFb0�4��+Z�`Mo�z2��ў��"�[FB�����pϾmJ���ͦ0���y�ݦ�&x�QMHW�#ڴ*����%���{�jwz�xa��8�2B�J9��iY<[�I�E��eo���׍0��)f�����G_[��p�����=�C�KY���fa�@n7�̓�[������5duZ��8��=�P.>>��tA&Fp@��hBR��͚��)��{b������.���r��s?Kď����j��KlΞDKX���n�,)n~��h�������f�~�4\7���p*M5aQy�̾���(�{8�w�\�_A#�����i����s�x�w��h��G�ɨ�n�9���k�-�Ѳ.��E�o@�Ǝy��_�~���.fT��;��3
c�d��^�Z��`&���8�j&'�8��?�b�w��Y����<g������pl��U�Q�|L�F��۪�<�FT�yJ�I���ә��9�i#�H|�����9_$���9Q�g��a4����è{�����	��Ui��O�P��������XIz�d�+�bV��h�b�t��?>�~*����^�e����(_��+�h8T�h"y��xK����4{Ȅ����ݞV��cO���K������fW��ݫ�
V�M������u�ڷZ���6�>t7yB\1G�6�^;z��d�Ơ����jό��k��?���>�}$�$�['a�������)�����|0^i�49�/[!�+�^��ϣ��*�_�������?(�����5(�[��5�c��ݘ���tǵڪ���>�W��ק���[�(u=�����$���+|�K�&�2��3��PL4�P�%��/�V�q]�VpP�
�.�N3�v���"�
}���AH>8j����9P!)vpN��,��ƿ
�?v�H^Y6y=z�Q�����"����lh�����ߍI������u��ް�n#�S:���Ʀ�ݿ�UNOMmx�����IӲ��8�	`͐M�[�rP5	�KG9��l��D��ʮ��倄����m�צ�Z�1���3GD����Z�4�g���dl�񈵃p"��ȣ�>]�K~��w799��v=^����f���e��B����M�SԷΡ�z<~�Y�ڇ�~:1����h[���4.�ƥ[^ة�׬f�����~�$�@�V5���S:0>K�+��o�W�UR	�X?\:ߩ�{q����tb{�D���C�T*Z�k]��5a��>��=I��oo>��� `�[T�F�j4�J&X�l2{��|�U�?A}'�g��Yo�|}r*~:7E��/�%����v�#ܝ�Od�N�h�_�����]|��s
صV�[����+���̶�*D����Uv�2�/�TQዿ����?� �����M�BF���kXsր����F�t��,fV���� �r�'6��=�Mq�4m�*�Ie����jܲ��v`��A����?KwY��}�C��H��Z�?��'p%~{w�u{m-��^�]�Od�|g;-�K�X]K%��o1OJh��'��D?KfD��i�|E��v͡Dua��=��%_~21oԾ��3������RF�Kxv?-Q/�&���f�r ��Mml]�cM,��f}�E�t	�ǋ�d9Q�����Ge셍)邾��fR�~�or��WU��PN>��^�Qc~�	���Rp�J����Ȃ��չ�w���m3�+1�����$��6W����G9�0��ps�*���-�O��Tڿř�*�;�ɳ��P�p�����:L��J�v����_���C���}yPh	��]�k*+*$�����\g:������4��p��>�R1w��M���(--�w2���%/ˇ�ձ�F勨�s����g;a9i�7�/W��~u�߯;b{L��g`��������f94�ż+[�,�cV���5A��1�⸕n������~��>�	Lh�,�VL�}��w�3���S�C��~�rO��r���pt�j��'<3Tӈ:��;}ۤ�A�,x(rf����?������h(ֈ�9�ݏk�v��o�5d���/	 ���ƖsK%��K��^M�B���+���[2��Y5倬����e�[�'a��"@��>�G��Lnmw��;Wr���tE�EvMZ��NK��N���@�8ua���
�%}^��r]*vݗ!i	
�ا^!<��K5eש�elݦ��S1^�gK�����<>�n��.����>Yӳq�����ַBb��j֤�TM!{ٲjZ�]H�v=��{q_�893D�[>o���+��p� �����pgraoq����+M#��|֥y�`�o�g�Ƥ�9?���.� ��~\L�O������������}쮑v��C�h�U�U]^!�����כ+��Һˋ��M�È9^V�e��P�ޥA)�4�S33boMס�ź��i?�?�=��7EP����K[�Q�o6`�Ӕ ~��L���U �4f��������)G�˯=.�y�7-�s��g��)i�}�;��S�Hp�DЛ�Ϳ!�k���N�u�q+C���Ķ�ģ�ºK /ڷ�߼;o�'�E�q�Q� /�y3�3=$[
Yp1�07��_�>s;2qw?���S��Qs����׽��3��02#��<������\	�q�)�b�G�>�W�>��<�}����)�D��b��"����?j���|�R�����[�MPp�I^�8��u:�е�bqH.vk��k�]{��^�:�j�a����CE�m "�����e��I�����$�9�}0��`eޗ9�v�)����e����+�	�2ڡ���!��Ѭ)/�k�a�c|uN�����mt_�8�����ɬf��5dŎ{mc�w]��5�S�^!'��x:��5���򶿷͸�֛�QV�Tꢕҭ�z��U�������pb�R�\n��J�2��S�jY�Br��M�-/b��mmq�yS�Z4�<�g�3�o���c����o>7�'����N���"��%L��������r0�N�߷)�'���PSD�,;��<�}��M�D�Q�� p��z!�\m���z,ђ��DE�Լ�T�qw��/A	A�O	�N����S�e����5��Q�fZC��C���� ��������̡�b���B^8����;6�<�O��}�߾��
�����*��֎K��q��\)o��4O[^���aM�I߈!4l�d��0���M��뒬��0�dn'
��:�~��<��Fo`ob�L�|n�m(�c���̇@ �y;On�]׎2c�T��lt/fu����y]b�K�c��oj�� d�d��h��՟�`[`%�~���=Qi��N�J���QWW��l�z�C�6�D{$� �s��V�?�m�j�<z(��N�)l����)%*+�I��X����գwY�7ь3v;gX�C;�i(�ձdy�,�X!�X�	I^6i:7K���?��� ۖ]����VL7�.��c�p����̚�2.j��v��5ޙ_��~ �����J�k���6c�ZnFd�G @6uD���6�XMU����L�ܸ��|�^��XR	�z�-����� R8x)��b��08�&h��oVQE�Ǫ�><��PV�?�@D ��xMe�O�s�%&`={'؉�A9��䯘F�Úa?;::>An�x���:|��M#�%8]�z����zR��������R�ƣ>���V/���?,��\��w���⒙�~{\��KJ�*	���c�;q\qt=~�O�A���m i@��ZS�@�\� t�`�����}����ppr�Z�<��O��z"�~�I�I௭J#��[���~����a����dP��-r�ЭiS�VSB]s��U#y����111-�灞�2�ЌT�"�w�%ͤY<�(uS�{�աd��= [S?Kn_1����|Vm�>��6o��×JF5_N������{|6��aɨ	�Y��5g��W������W'q{Q\���m��:������2[w�	<(�Xz��
��*F�'|�n�agF�6�[.g����Ҿ=Q� J�eV�?r��Q�-�xnȘllo���i��ٗ��S��no�q�-�LԾ��I��u�����1���t���y��//��{��~��?^�y
���G�jc��s*�o,�;�\�4��
"��T(Ѡ��Ɍ��DF�ĺ%�wY޽��/5Қ!�1.��Ǣ�2�����2�?�B�g�A/��2�Br[��|h]��"�k��^&W]��vbc�ι��"� �TnM�����&>��XE�
��Ȍ3���nP|�_Lk(�zSA9J����R�}�&�1k���B�*�OW�-9���<�]��{۫<)�%WJba��u�2��_�j�C9��*B�ʠ�����a�������1���nՒ���� ��$��?���b%ڂ7/L�Ű�J�~�jO2K���ɱ�&���z�Cu�K�Vo#��vc�0[�dM�<`�d�N�::�]?w[)�DM��{�*u]�fW| znYd��i՟�J2�*7��%Qн�%�JI�r�S��o�/M}�zk��n�׻���s�g؄��a�
�'g]x6$黸�|Wq�tt|��r7��ё�]M#�5c�ޢ�[�x��Zȯ���nZ��b��z�*�]�������%]��&�Et<{,$<�E�JR2v�S�<�ɔ"��i�L䓏:o`�m��%��*�&B{����D���0?V����{���mԒ-��dmp`���H1G)�$0�0�i��n���;'+eݴ��@�7�v���x)��gk��P�L
f������Ϗtn�&ud#x�Q	Q'�NL������!��C�O�-Ӓ���� U�������]K'S���2�8; �3���OAn�I��Ro�H@���+\���'��	oJ�{q��)�^Ǚd��R�v��3���k��̺Rp��w�=� mu:%��:z����1�T�k8x�X��bюʁ�~K���I#O���: ��0�\�'#��z��J�v���Y��C�;᜗��G���SG�� 
+x�q{���y����u�3�`�Dy�w���d�N�t�?����a~��t���$\�jfi�a\��pP9*�j�P=�,vp�޽�	5h`s�o��l5�9���{.���.,����m ��Do�+�]�%UZ5=�/*ި�iN�*D}�>*-.|��� #��T AY���d�	g{�l��J�A������M��Y�K0�b�W����A�۞-%J���ďA}hI����񣨁oB9"�J�u�4I;s�7��Lhg���i���� 4���?��/<פ.��g�ߪ.!�>ې��ub��1A|�W	h�I��b	���K���,Wo������If�s��j]a��m���7_E���!|(�t@�>���[$���T�(uf�t��}����{�>�%��+$��/�ڵB�8�4���?i�8GO��3�Ӓ1Z�q�E��4��4��3�_%���C������5Gj���l�D��wP8<9ꂇ�,�[��2�3i� c�`���mO�{:�A�啛�$���4h�Z�J�Wh2gqJ��(Z�OR�#���zX������j�w��U_q�!���=��t�N��S�?�,�i��w[jR���/'|���'Dfч��#�`�S�u{ǵ7��N���[ެ���N	���q����a�����NOS���p��\�q�*�J��Ѹ|GT@����$��z.�y���_��*=��s>�(��E��o�g�b�o}�ƕ�̱�3�H�榦���I�#��wv�e�%)�̻�J�8@��_]�(�7������ڋ�_'�����ѐ���t����F`A.#�`F>l��i���6*B!��K�v�K���;~�>�y>Q�cc\��ې��.��`x1��K�[-�~�ȣ�c�~>�G�+���)G�����R��R⽈GE�O�ɑ@B�����o#��̌<� )���-����kk�t��$}Dx����.h9(lTxO�9t�yxxF��Ի��?b����#�^���u؉�V ��c�%��1^i{�ǈ�L���A���r0[�jE:S��r&�,m���oi��ͫ/<�o;���r�������m�L��%��͉����d�@�Ƈ��j�!@:�E�>�]���L3¿���@E�4*ȇY_��`�iJz}J�A����2���c�^j�:=��W�+۪]5S�t[P�5z[�.�y_�'D�]�EW�E�!)�H2����_�"�j�d1�e�����[f��Wf�^��s�T/<V�3��'������s��n@��I�U�#�f�x�D�����{�S`$x���]�t�?���4����#�.�ݏ�X�_ňX���^ g�Z`M�m<,�����/Uf-��K����F��Se�}]Hֳ��XޒZvS��K�b2E۽ٖ��>I�B�4T|�O�_Y4�#�Fb��%v��>
j`n��_�ǀ�Ԇ^l��l�8裬����m,M��̈�87uJ��v/�=#/O�~5e?��QX<�nhږ���*R���ڤsg�]�;��9��A��~=��W�����%|��;`�9AA��Ę
!fڋ�p`l9�jTS���+}�#d��6�`���ЖL|�|���-��"��l���_L��Q�T��$��ˎ��TZ	�Q>Ŀ��x)�)�UTt�[��E�U�Mh�N;|�� V�s�4�&m���Y[��4u�.������h�U�	R5��97b%i���8���r�MIIy��vh~6����݆��HA��R�0I=����kc�VGQ˙���۔p+
<OOO��Kb	�~���
 |"���q��bp�����5~�	ЙK�z��V[AE����#�:�n�׌a�oc3�8����V�%��s��d�:���-
�}�ֆ��!��e&ژ��>�����3�sЧ�����8�-����(Y����ym��^u���fkt��Lf�?�XQ���k �~.�иƃ-�t��4"���\��6D-<^�Cs�Rs>M��h?�0�G�!V�Y��n�	�$�F9@�@p��6M �V+��?��~�o �*V�@�����g��J(ӴV�P����ػ
*�p~��]קގ��j����m^9Wֹ��{ƦJ^-ܖ��9���O�э��#� ~�l��KӦg6�{>=Qs�Ư���e)H��#O��p"�5�Tlђ�硴k�kj�#5Z��v^��8��6�MS�����7�!v�Gn��j�W]1m܆��&����d�&���"*��J�b���&8�i��A�t~�⦺�/_޷lj����o	R���Y���T��u<(�sy	��Y�Q�}�)X6�A�X�����,A%�AK�Ҋ�Htl���L�!�
iB��H�B��e�_�����Ҳ�9�ڽQ9��e��l����3�<TQ���8�&y̦��}W�" @H�ٓ�>NW�|u���x�K)�s	�����y᫏�� ?��E�W�<�pKħQE����Lo��?�g�Z��A~��S��'�%�W͢���ݚX��~ �(�M|"�1�N�i���,�����<����I��%-�|cJ[[�|B�<�^[1D���/߿_P� 	��m�'����W��e	�FG���P��^��>�,�:f��i^@�@�-�J����;��k���N�N�F�y����ϭת��Z�Q��MC�"�+G���ZC�ԇxa�.$ߓٙ����sߋ��1�������GK�yt�2x�X��;</@�icٷ��%�l�--���xo��1�Ƈ��jZIQ�?��9����7ʥ�&�\s@�@~x�~�^� �r��ʔz}���qW��K?F��=�)���+�X�K�Я7Yެ�x2�C�[ٟ>-/�Y����>�vm�L|~�v��~WcVSS+_m9���_���1_׍�$ʓ�]���OF'L�X�j�۳k��ު����T�������+ jCCx
�ʥ��X%⮽1f�0�@Ĕ\�[�܊����.�B���++�U��u���F�z��Z#?@�hT��;�8�>#e�)#�}�R�[�I_�si��/����K��Q~��]4�n�ǰ�n����ڷ�=b&tU�NM����&��-˱����fK�g�gj�T��Ѯ��2d�T���o#Tݨ�\���	��A�R�ٔ)�����/3�g��"$  �������.��z��RQs�Һ(Xb~�p���]wW-/��a>�ͨ����3���(�I�l�ǈΥ����3��z�f:??�˓�}��3��A����;4���L�p8-����D#����)������~KN����Eo����	�~�uW)�Z�1�kc����y :GFn���b����W�ڈ���f!��8�0��q�k� ����w]_o���X�Ue�z��ӧ���(���P$��t��,7bRŻ�]���6x��#�6�������p��kq/���U���62��!P!?F��~��vWu�[w��G������qq�j8�#\�ש���,%�����|m�*��o!�$
H%�n�e�ОhZC�`������f�J)�G��FQ��j��S8Sғ�W�3,8b;�A��n>��q��[!0�ae{0Cj~}$/�V���0��־���=�? L�&�)�.}5���bi�u� ��o:�����;YHV�
����h5���p&�:f�b�ϧT�,//󤕗Ӗx� ���dg�$s�	���c��ו,�
�,P�h��4T��Y1�)��L����������eI��j�dw��T/ώad�%��r�7q~N��{V
M�t���Gg��C�z|�Ͱ�n~mm�2��DK"����)�dP�-��!%�����.���xv��A�SA����'��p��2*GlW�Yw�����H�����Ϛڱ�庻�g�,�֌A?M��'��Ƣ ��)�纨(�3Ia_%A�q�|*�KM��&!h��t��k<�!�Ȫ��~����D��ϸT�y���:ؚ�٥��}�٣���*6�܇�t4$�!~�#�	�7o� �Z�t����z�����k�ð�/�>9Їz�i��"XK��8g�����hfb�������Erɜ�uݤv��u�3�@������k��@B�-MB����ʜ���%w�Q���/h:����yx�MT�X��|�|���R����<��[��sr���C�C�+�dXXlfd��ڎ'��[�|�*��X���7t6���yBrrrU��5�V��iq�l����.�`���y�PO��E��Bu���",&������>Sh�Fp���m+þ�=�o��.N6$nEx�	��q^;��� =���@�U��-M�P�����������J������3��t����6�JO$��ԡZ���͉RWg��&��>^h��d�Jff�wˬ q��]�9��s��5��m�Տ��Q.�;a��F{}��_������O���V�P!���n�����nX�d�F��^c5�|�dGT�N}D0�'��1h5<ߨb�>�w�aS���l���ɵ
�
5�Bp[�_@�I�.����������,ٓH��{k|���zbF�mkkk%��7x�S��Ȋ"<��C��sØ��v���s�<�ڜ�x��:�蚙�Ԑ�&�y�H���'�W �Q��h��C���8)R}�3;��u���D�)BY��a�'��h�-,�T�?��]A��~�$F9{��I�S��v�ZH��� d;�U(\-6�*�5�3����P�QX��&�IV��@�|���~���x��{#��ʯV�%Ȋ�����e��]�g��G$�;t�� ���s��cR��g����%T�;������JȦ���:��"�/�u5�iֹ=��c��h�g�3Y�	�}]S���}(-'g�okrO��/�>�)q��-� �!=�^D4�	��c6����n��� �>����!5\j��Sr��O�eP�v���6#o��R��7&zlpP�q�p�8m8
sHH͆`a���"�֖W����a��v�7@gi�-�k¢ȊuvK���5���Ʃ1�66�sXϷݍ�K���k9��^���K6���{ ^�Mq�6___��g����{.Pw����R���ђjL,,�U7
N~~-��a^��_�W�g�W�תq�w&)?�e��pv'���"=�y�j���@/��r_#��\���zA��jX�ܧ �
�J{4�ՔƗ"����:��?g;ڼ~t/�&�o�

J�-�)�<�sp(����*����R�#r�������}GTT��P�+�ט��@�7**��hC�y�^=,��xcw���-
�K8���vsK=�/ƹC��߈m{��_P�_�e1�|�˴WC�4Yu��43�7��Tn�)�}Ң<9ԘB��>�ߟ�@�h9�\^���\���l���t�N��@�7ǝr�h��s�� BR�CZ5�o�cL�)��;�F�l"��5����<�6G�Ź9]���voo��>x(9�E*�����.�Y��XS�56^>4��N�pf���^^�9"�c�\����.2����"���i��f��ˈ�|u����t).Y���	uO��1	���ɑI���C)��c9��1���ɘn���Xﱽ�Z��g�Jo|��Ch����O������:���׌����T�6$x�9�����l�"�j�G�cc���r�?;��tb^1�D�
��k�"M7��V)���>���.+��G��WB�S�5���� ��Z��	���]��j&��-[�F5�1�$��Yz,�������t�!&PbW����6Z3v9[�޲"pX]���]�>�mr�ňhA�C9u��k	�/4`�;���}�Rp��]0�q�*g	�,+Кz�6��<�ei���ӕ�M�I�rcjΈC����d=τ����Ǐ���M�S���r@8WV���vo ��aghh�T�45���E�G'��m7����n+b�$^�*��3$^�<�52r���p��\�"� V���j�1�]���bu���LzNM��{���v�,�I��^^Y������9�]�Br��u5��,r����n��&c�@`6ߎPǶD�:��h���I�a���N3���˳2�D� �B��gC��7-�k!R[5H���������-p�^��M'�4n�-�Q�ȒӢ@���u� ��&�j:���G]2�Ai��|DX��p���)��K�#��KL�Q�־�ug��q�����:�i�1-*�"���F^�q_8_� ��Q���~��t�=�?Ԙ���q>����ё����~p�@k�ޓk���,c��K�>����B�ƕ�:�rb_&�G��o����e1Io�<j�r��3�IȢ}Ǧv��_���_�޽D(� !����VS�4��j�)��j�g�*��a��K�7j7�OHη׶����㓒�TB���+mt:ކX^;��	�.X�=�D �u�zw��)��yh^ޫS�t��_@)^�>*"��p��b�����0AX�%�k���!��2,�5�y扖�ix EE����Ga�eY![�+�P�C����v�J$���&�O�cӀc���o�����'����}ٺ�`4��;�dڇ��v��x�F�� �x���a�L�k~�<-��O�4��J��7|0~��z�r5^jmP�|[ry�]�S�6,�~ߴ�\�9Z{E��|�2E��d(kzĽ��q���x�� }���t�N���^*H�W�DLB�^��e���p.I9D]�;f�E�=!Y���^./�{�܅��'^*jzz�ң��{PH� ��b�ŔA����N�d �������N-uH�u~�]�S�����:MG�i�N�{	"�T��%X8_�v�v+(����K~p���y��l�l�;��mr��p���Q�����̭�V����8����㇏����Ŏ�is�����m�YL7�K�y��¸^���FՃ+W��?z�?�7��<=�>8nW�$y�	�+ڜ��������}���)���ߞ�i��/kU�Z��yo,����iV�k�}��p���y/�N?t���悷��G�%�=�o�f�n����{��/.3#%��}�P`�+4�������y��dKv�������\sg�.}����w�z!����YW�<y����\���U�{��~ϧ�ǯ�KCh� +Z`fק��K��̎<�z�ҥW��7h C~랸z���2�Aj������g�7���s��-��;o������]�qήȣ&34.a�uK.�:M�y��������a�]���]���������w���Zs��!??Ƽyq�9�l�=�
s�5��m˛;�Y��q�̙����f������/o���goZ0#L ��<�����{��cv���]���9���e����L�<NR��d��`Q�9��u�e��m����2L�9�������Ƴu�j?���?{vu�Y;}P.sQh;�����w���W��ŋ�a��~~q��}~����d��h5Ao�� �]�������f��(��7m����^��5�O����'[����d��+���"���_�N��?��9�kkj�|�7o�������<�����i�S�4.M�e./%�%����tFU��m1�����?���#fOR8|y��
���8�0���[*�{0��o��5����~�ž;~����C��!vF@
����<٭�bRa⁗��O�8�ߢ�D�ךf"!�ǖ-_n�<�W�
�΀���}�z=��[	��E륤��nݿ���,a`cg��H���q�&mt�FKÂN>�J W�4=zԾO�m��,`�������xm�t��mѓ�����j��(xsc�6;�L�N[|��5�9f����ۖ�
)�����VvG� uȧ�	�(P�[�q��ՙ&R���������N�g!wz���B������p;����yo޾�����_���=����#P������ւ"�=y����{��N,*��Sbч�����|�V_�ni}%���G6��/y�Ƃ-������Q����>~���I9X$��b	��J�r�dVY�cyZ*��������������ރ��&�{V����߻>�4�j�������}]߿��{���p�~�8��.�r�.��߲���J�j=���s��^�����f����w�GYw�_�w�v��w�q���Th���L�+L��˥���J)��OO�k�$v)����'k�������gA{�Y	�)��w' e��$df��:��3��8�R5��d,2��&R�U�>!�n�l<zvރ
b��(?���j�lʴ1�.\�p�L�bM�h0ˋ]��cEρ�T�$2��΋��2��v"���Y��T6]q#�\��& ���l!���������+�͍�����/qJ�̛��.Mf����ѕ�����Z����L%�T1�sʀ9�g%���F'+�Q�yw�B!�X0OeN���'�,M��ߩ?��V��	߉_�A�1!���y��z�Cäig�����:`4��&�A�L���9��Y���3�����e�SB PK   u�KU�b��� L� /   images/db75ecfa-5437-4ae2-b047-1b58b40ff187.png̺�7�o�7;v���F�j�ثfi����{EQ{�&Ԫ�6E�E��B�(mS5�(j����|���}��OxNN�}�+�\�}�z�_#I��]z  @��w�  � H)��đ�#��@׳
  ho��$���+�{�B�w.�]��s%�U�u9#�oIIIKI��Q��;��WW�X
��L�%��q~﬜Ӳ zl��q�:�{���������/�־
�c�s!M�,H��_?.19^�jz/7k��Zl:���^v��>]w1.�_#}]{d������*6�$g���3n�9 ��+$D2b#cz��Ҡ�ޤmUu���{(�������+]���S��=�/Rm�O��vx������h:�a���x��;I��r� �$��Б�1�bZ���B���f��7�b�՛n�^�#`����P\ 1q��]��W�C��1ܖ�dc��� ��J5�w�k��c�6h�E�'6D���b(s{���M��W�U۾hz�7�V��36Fdv��F&��.�m>����Mg6�\Ԋ$�/;><H�Mi�	���|mJc-҉����nU#
V���q�A�%��'zNN~/������ �@�j�(ɳ2����hl���)T]�bJ�4����׭�ky�|���W�x�}��e�٨�H�h���t.�ȗ'�PoQ�6sT�'�M��4��������{�{X���O!�AS�C�u��O}aT��
=
U�Z
i�=i�}NR@G��Fd;��r�d����o�P�Or�!Nt"'��"���ٯ���Y����ؠ����ƉS���.�!�$uo4�g�͆۲jN�?�l�X�Ւ��x��fmY�DV�Q�h�����W��Dx\3����m��j˕P��<b��#j� �ؑ�ȟ�gK�`|Ť~A� ��η���/�:A�3n�Y^ )�� �9ج��3	����WF/��$<���Zc��l+��x�EX0]Z4D�9"qC�a�X�W�����L�Iѻ�#�m���Tչ*���|(V
<�
1���n��phᜲ�Lh�����Ӎ�2��1\���n�$�Z"
B�|@�Qu��f	*���������W�� l,�tD���}��""|��1�]��M<7�nt6z]��N˓lX�:�X2#��x2.�X4�� KVJ���T�r"j{�C��f8�oƀ mN��ƿ}cU�j��ذ� G�y����0�z�Em���W�1��\5mF�����䍜��C�{9۰��P�
��-Ԁ0$���>��MĶ&Y����o���>W~pY ����Yu1�X{@��?��q!Bq�?lͪ{�dǑ���R5CPT̵m���xaѧ�~a�`����i�R鑧�N�v!W�����ru��w`��G3�K��}�������M�M;#�]��gS��.{{	�+��.nS�`�ip4qM"㔎�Nu��o�j�<"����qQt�i]�������.�W`h�Ǥ��ן�����7�H��ׄS�����upA1��E^�-Y+`51�tƦqсJ`7����@g�m3Y��Pp����	J�)p��:��t{��u/��n�w�������!v���W�u�u�:Z���h�����>�O�;+�^�k�y�0Ȭ9@��o�G�2����%1�h�C#yb17�7&�__�\#��`b��OY��Fn���:�A/�),xe�RF�A�l��4xLξ6�Q{`p�K��u-�e�q%1��NݻP������!����ؘ�}>�`�O@���s��d���u(����J�X @�UJ�ֿB�N)��߯V_&:�]s ����b5^��M�����ݓ^p�r����V��8��,�l�%��ϳ2%�����3�X	ޝ.Ro0b��wP�ț��
�������Ib ]����l�bI�O���dѦ�R�s�TIi�1��_��]z�0�׵=M8��n/��]E��J�B�h��=B���缠�������cX�����}��s���54������ ��H=��J!��oi�X1�&����U"�
��(���(��q�#�20��(�w�%�N}W"��&U��#f�+Z��Sh�� ��ߵUSQ����bZ����"�	{	/�S+*�L��"�l53�Lʓ
0�,�[��h��� :��<��_j%/r�D�����n��yƽ�������O>39r�s��t��W;0�~�Ո�e���%$xηk��Y�s�5�o+�K�gSl�'��4W��5�N����rZK��O��M�B��(��Vdю���|(��G���֣�`��� ��%�H�]��6p� �]ɆI�o}Zs! �oy(��:�A8U	�$���_��rߢD�/�q�o$�o�LI�� ��]H�����%K� ��w�ٹ8	��	�0�g�{�;f��w[Jt�M\�^�tQ8,JmB��	^h���x�꼯��"u #S�CQ��I
�j��]����RB�x�o�w��]0|Ո\����� [�!u��x۷��P�����\�8J����i#����u����́��Jo���y/�� ^��7�M �^Ԃ]J���(87h��{���P� 4{�P��5�6�4�7������YoG���%�	�3l�13gl͒9lV_?���=6�g�=�o�e���.� �� [��7�f�mq�q<�s��Q��G������h�UM#�#�[��������˗/1M�L����E��������v��@�O�~U�*)j� +Aَ}���:f�8���F'Kr
M������\��������;�F�yq�
�k����� BH
�(�W���&l�t��V1�1{�p��uft�A��(E�`x�'LGb�g�-w��.. ��/�r;Ft�i�c��
Pc�+wS�s?=��*�թ�7�� Ւ��z�L��lU�_�%�\3�	����?^��CBb�AF	���wH��E����,+�F�n^��=p�y���K�������!$��ë������Ū�2���w)��e$�0�ܺ���YFmّ�u-�F�Yl�	Jl�\|f蠁�w)l�)8F�b�.|�����h:�x�]DW��L���t"{��f˄i�M"�*�#K��A��\�	Ʀ�<����y�DY\Ht k�'�3��v�uA�U��W�0��&SG��	�NT����@u�PV��:E��Df�]z��^���2S\Vio��l��F��z���-�p��� ��P�Ts����� s�++�J:�R>�1��ܐ�����ľ��$�Q`��$�j �ʪ�J����qa��k��%F��m� �)ʍ?�]�V�&��\xu4͸y�`*:n^W�L$������Q��4H�<�`�/n��|����*>���/�bs�/r�)T�1^� ��G%I? �����}�w�V�{v����N�7�����
�	��z�J�m�S�\sW8�M�����H�C�]����
�D���}����I�hwHق�@��?9�ߟ��:��S��tK����B<a6���E�?1��g�K�Ř2-��ܫ�$�>�d3���	t��ҼU�h��6.H�� �?ʌ������5��߾��1�ǝY]��kX�q�3�������3��(� h_��n+dO�ǹ�	����p��:)�ta �N�f�5M@���}�
e/g�u[ݫz7�.��	sGx���yS[;�H�m'J�]�#PM�"��:������FzIz�Y9����[t�p	bV!"v0+:�;\�p$�s���xI߷s�[_��E3�[�%��ZĻ��=�h�!�ݫ����˲�8�Vh;��� }�O��jK��x���Ef�+���b\}-��K�uaw�M~�,�!�N�wI���8}q���;z!�#����)�?]�񼡂dA��&bdF�H���歾�y�8=B�������6�b�1����U!��[r�N�ç���,��YV(?��ˍ,�Z1�<��et�9q
w���#��gf��'��ɠ��z�F��FfN�s�0_�2������e$ֿ�B"�ݧ�a:�b���<�z�ݓ����$S�K��h|�,�X֦z5�v1D$��ҩ�և��j�������Rv=�`qИe��ab��� [􁅀�����-Ϙ�������~Qv��Q��E'�:&^���	��^'��T����^��v��2�pST�>���{(t��%v:i��o-��û� �N�[��2qZ}OQ��G:���I���~dY�(��rgȣ����}���>W	Rt�� B_�
f���ƈu"u�RmR�h����W��|���� t�F��	�z����,�p��{�bv+�e{��7Kn�R���9�1O�	202��j�����~���?B���4cgWi�U[!�!+c�EH\@qq�c����݄�Y4Nn�������ޓ���%��\�X0+a܉Q�%B�3/u\Ƥ�!P����G�%A��o�KK�Ӳ��r�a��2w.�{e`���97䥙����Iv��-4g�) nV�&�ަ�C@Z�����,HKV����z�}E�`gt�M砶�\�ds��Uq,�w	*,]˛�1 ,n(�LV��(�����?�as:(^�*�r�V&�/̶�����0��]N��"3��6~�G�n��kI���J�Ԇ�544�*b�oa���Hz	f�=�!��ZX�,2��mK�B���i�(_^�U�
dT�V*?yl���4ǎ����������l�U��LK�1ng�>D/\�I/?F*HmY��<�MZE>�1��k�4T�b��l��U����+���?2�'�����H}7������FԞ����/�>����-��G���1a��{2��/7�o�:��+em��.�p�=��s�X�]܆)�XT�1�i��]���^���AT�?}�7��]�
��ׯ������=��L)ѫ#��3�t�D�r�A�"�1�`$�FdFx�y�'9m�؄[�X��u�@MF�]$��;V�G>}��܂ $���2jg�.��>������#�y�dJ�0�mIr��n6mu`,��lv�XN�?2�(Q�B�x�Y�&����W`����9�|P}���R~C�J��<�V�D��$f�X�+Be�?�Q�` �,���'���^DD�=�@��#�7�ԉ���֪7͖;��қ�w�LX��H�W5ԟ��,e�rRz� ��ܟ+���8[���|Χ�o�?X�U�X������\ۡ�������G޴Z�<��>��Y���<V��W��� �,I��Ⱦu�`r^�X��/֘r��D>Q��'���gs��(�����'�>g'+x���CS&!�L��-��CCZ;ϕ��:�qn�����Zp������q
� �S��d�-�Բ%2mui���`0u[��_�%��ip=QF�*N�-�X!����1��}�Xq�-bN��QN`��Ǥ�Z�)2�[�q�G`nii�ˤ���^�ꇗ����W��!�V�0��J4�	480}�y���[�5A��I|C@�r ����j�@Uת�O�U�YG%������d.R��Zz�
ISM/�F=>&���r������%��h�1�~mq�œ��9)/�:��^�pR�����eU-)�C���gO�����o2DtEb3���-�C�.~��]��.�f�[����k�Bi	W�tp,�}�+owͨv}��֭[q��r���+cL�Y��?��I�P[��}��y�s/���1/�V�G��I|4}�r!�C^���k�6�h���?ey#Ę��>�k�;n��h^���rIE� ��H�ɹq��Q0U7zX����w�7�O�:!����8����������F�YB���ON��x}ϳ'�;s�)�����}Jf'I;Ѝ�&�d�[o�l�T���n��h�	9��"2�g}��P�����]	�k��&��dB9��Z�IԖ�*v�[1t jj|�r�6�)H�x��a�핓���`��������ԯǑ!5<=K��2^V��)��c=�h������	d��Ox��{� $�-d/�tg��WZZ8C��g)9Г5�d�9�C���<�
���-�T/���0I�M�� q�q�>���EeV@
�^ D�˞��T��N����`Mq΃�(/3.�{�=c�ga+@������7Ʉ�/ �Y:�MP����(��(���G�!)�7�6���3�{e��pm-���.L'�w�< D���z��ǔ� �u	����9I_m��lĉ9nO�3���l@Y��;W��|�fÌ��H����e�--��_�ѲP\�c�����t�BL�Zv]����fYuO�.i�2@�Be�����a|н;���)0}ô��&$Y���c��.��g80i��Կ�&�><����W�s�L���Ō����1o�ވ���]'7�2ؼ��#�����l�8�zIn�S���}ݟ��o��_-���H��ߖ��ڸ�v�%�g���,N21��~��h>��ir�<��㯂�O����?�=𷹅;PWf2=D�,�s�V�����H6 XK˂�������wl,y1�κ��O�ҳ�m�Z��B�cΤ� bn������<�&��rp��_�)[�^�������K$���`�$T����J�{a�md��y��Pf�HI�n^Uȉ�w?t~���������gӢ��L(8���+��O?Q�j�9=/��^��x
4?����/^Jh��^�w�����W����lu�-�ݮ�<c��F�=F�-�C��(u]!u1��g��x�=�b|��4�*�|��be�����CV�a�����#�p�w�>�{�Ef�&�d�Ͱ�RM��B���7M޺dBS�Vg����E�%ӱE^�L�$D	�Ư���:�ؾ��Ô���XS�#f��wg����1��f�3�����O�͙���9��+�ݠk&n��;I���� �}��+'�O\�/����Re��<:Hfcuq�\�
7[�
=/�7X&�i�CԬ/��F�|���ҳ���}�:��8�(<�ŲK�:�_[��?��z>2%�� �v��N�{��k�������7'I��DF����1���c��{�%��pP"�񔔟�i���`���������	�bE�VM�ە�岸�y^ ��^�0�puۢ�T�v�C�E���ל�+
1j+�8�_�=��#��85W�s�)�@�c�_:��N$U�ڟ�~����`�ؖ�KWζ����0��"N�^	$�۰$�}n�����7� 7k�b����Wxi���9?�s���J#߾�vH0f� ���� 1X�CΏ�0���kL�U �vʜw��󌴴 �7�6vD]�`�-.��fM�c�W�ؖ]��s�;�L�GQ��"-:dH��yι��C���"�s��Y�7�0,��wj�ߔ1V ��>;��ZS�<3r�
J��,+2���[X��4�������'%f�j,3Z�:,.R'�!��L���%{��ʇ��F�r_���� &u�Yry_v�D���!'<�k�Í[���A���@���xw���؍MV��X(ݮ�65�V�������sI��e�*�\�&0���c���|QN}����9����D�Jv~4��������'�ɛU-��R�b?�C�BY �J�,&J�l\�7�[��.[ad�{dn���=���`�]�1���cF�r~#H+Lh�״\~�c5�t��~
�	6e|[�=澁�7���V�j�ϫ�B��G�H�5����M�)��^]m&ʝ�Ex�0���!6L[~�qWQ��e(z5�|Cv�]�m:JW��_���:�^�>�9\����D��gN�����ЦK
�;Z]��8���n�lk�~���t0�1������mv�������j�=;V��U)�gK\	��TU���Z��� ���
�� hb���Vp��}��MW77����&�
-e ���M�`����<LIi��ؼ���d�i�a�{!M���B������iM�g4KU5�m!���<x�rsjj�r4`��v�vJ{��sŔZ��%���e��n���3�#���1�/�#���9����o�h�%Rzg����м�+�P��YN�u����&��*��n&�ɚBUl)��~F��Ԉ7>m���Lm���+>���[���)�tS��tY�G� �!9`~>�n����Н��㥱����W����vA��¿*|����j������$s�7ԧ{Ml�b�����dfx�x�]ْϕt|k�Ͽ+Y���4Ȗ�r�%6��6B�G�L0����S_�S�Ֆ����1 {�0�btLw��Tރ��1p�M��Bx<�oANtrɿq�C��"����c��iퟫ��ў�f�_�N/y�L:��4�}�T���Z��!�n/6�tܻ-|cy׍zc��bhq���9�Ad�
��D���?��y��Q����;�Nӫ��۵�j��@�D�Ba���Pc�f�~���kJ����o��8B�Q�����g��U���G��x��N�	4y�MV�I�7��oHG�|b�&[^�t�ru����X�eVִ���9*02iQ�O3/g���Ȕh��p%� �P�~��s��/�	�l@.X!���^4�Z��7 �2ٲ ���Z�E_����O߶ή9��������pf�@�R����M�ψ!�����ɾ+�?d�.V��kDPM��'^��MҶ*��Z��Vԋ+��ʄ_�)�!���]����XA��X�6]�L3��<�]Ol�{�=�=����F����b?9�xIv9�[���dJ��w��,]uF~��	]���2���r�����?t�>��T{�������Y��r�b�I��3��"My�;�%�p��)&����{(W���� 	_�3���Q��ڡ�1wg	j�����H"��|��<��[�D��Y��T*u唩�LdF������/�g�w^R�"�l �f�z�-��Xd1�����@�;5mo���ڿ�iD����y�8��<7j$O��8ӎ��JJ>�x'�*���E��1B膢�=a� .,寁��C�����
���F:���ʝ�cmqq������p�;Ax��vq�$N�!��*[��?���p�s1I��Q����-���e �1�:��dTk��y	m�Wݷ_�{��y�"� t�{�x������~�V@*0�x�&��Q}����O_��n�-<N�m�(U����B�����` پ��X9�.1u|~����t��RS-5���?z���]�K!�	^bY�2��ػ��w,����l�:Zߝ�O���x�8�U#��~�I�4K@e�c�g!\�� #�J����bv�|B%�U�l)�a�/&�ˣ��#���j�)�A��c���'�
��(j�ˌeSGyd{Zhɓ4���Hm�#�Ә��,x�=z�.]��{2�o����=qm��SR�����C��,.�x��=��r<F�1�J�����@0��`�~s?�����Yggf�Θ�������Z�Mɚ�`�=7kWI*�
~&�Ά�a�l�)��M8�v�EEb�p�}琸��lF���@�=��9(���@0�A=����l6�����sK/߳�K4�O�I�s�##>n�on��u�*��lx�H�_,�4�T����$�4�|�]�)��_�F9$�,0�u|���vΕ����F *�J���Kq{���B����{��̓�~n}���?�3�����bޖ%)���z��3��*��v_d�sj�|�i���UD�.|�ٮ���Tk�h�g�K�dx y3���>s��� �FQ�MX�pOB���(u�?�qԪ��8O��,�t9�d�q�S�H^�+ߎ��/�� zQ#�꽧����%�S*��Z�VC��5����ݶ������,�.�0Q�V�,�=���������e:w7^��Eo�m�;K�� ��=*�<��:���J�ܩ�{��F��WqOx|�0�����A�� ��ٮD��.	-����0fb����_r��s܆~5��0�I���9�]���������5ƻ�Jր��pIy�x嶹w46"�mY�;R[�(���u�nC��3�����߫N,r � �s��n~j�l��U��H�Q�$`u���}����x�s�ӽ����D*-]��}:!t�H�t
f��zXc��
��ދXߥy��XQ��$-��Ć�j�L*�M�V��3�S���� ��Ȍ�7>�r���m�y��GP&˂}
�eV���\]��k�����'��&~ 2@����������O��8]c�0���¦��M�3��a�dĔGe��]׺���|=	w�,��g��,���Y[��ϧ4\*K{�{}�B��;=�F'�t�g��;=��;SJ��@P��oKQ��?m>~\_�|]��Wx7� '�y^�(A��=^��#�S���0�'�!�}�c^:���̹�T��,�sj��	@�>O#f=���.L�|�*#o�,�;���n.��0��<,U�^~�s���Npd�mFk�4��{�#��C�}+!�[�yЛE߇i��e?WܻK��݌�X˃�����N�F�I+�ܽ{%�����I#	^Zj2���o3�K���8W;.���w}|m�k{��'kX����HJ/(�OH?����2�K|���k�l\�D�������0��66��,�}�a<�����R����Ȫ��ߓ�3*�_)LsO�#�}Q�^N�"�SXv�U1��N��P�<*��oY8��*�ݾ�ꉒN!��t�
�Dn��F�p@�m�I#���;���,]�Q��4a��o�$yY6��``���^.��R�s�y<�
I�Z��b�-0%��a�A��׿m��Bt�"1�E3��6���e�c���_y���Τ�2k�+���ˠ�U�A��q���r$��B0��M�cW���Qۍ�sǑ2AN�����AY����"䕙5�T	�w��4���t��9��%�# "�+�I4���W'�B��7ↂTԑ�tIJ$3QO6��h���?JJr�<��+c��_��> �I	��
k~[�i��5�O��{JS���FC2c�4��߆/���^��ʟS�2?
Vذ�� RM�N��Q~��*�t���vQ�XG�F�}P�Aɽ���I����+�>I�4�����[-I���[6\����^�	��j��9�;���w�_��/*M�3�ۺ~�k��v���l=���c�?����.�����o��o����$d���G�=���W{��{��ǶM/&׿��<�ƪ|�DQ��+ �������Q��43k3t��C����g�i}h
�N�o����	���)'e#�����p��`6:�qu�O�5
�M��2Hu����7q,�nvLv���yv�b����WYJ�v�g�����������p�F��9Uoj0�C���Z���a��RCL0 �f���5��	��q�d䂆��G:�4�*���l�" �?c���%���u����[͡�q���a��H���|�Z�
�P���A��V}�F6���I�_�QE�}������؝�^��4[���E���w��|�/XR�)k��A �(�A�����o���	Zm���T������ث�.օ�Y��a�ћ�������#ΑudK;�wK�x+/&�X*��©���[]�]��_���3b"	�8�Mi�73	�	2.��N,׼Q�%���ط�޷�^l��L\� R���K��čN���.�r�5�Oo��N���W�AX됔�-}�V��Q�� H�Z��hv��bk*�=�lrdN~��F��b�v���7�hM~�^_��F�dd�[Qf�I���$�;�&��Ǽ"��E\K��)�t�ȌE�#N\��Ii`��b0�vG.�s<�G8�n����;����2�M+��:Лf���[{�۝��h����&�|@}���v�ݸiX�`>�����a�HZWpf���æW��#�*U���U(�w:K����E7H��痕	[����R���l��ops��s�5=���ۖ
S�BP���/,u�A�`�Z�ƛg(-�<cS�)S�x��.D�y�Og������#�6��|��1�����`K�Yr/��z�Qׅ���c�+��E��5���677�R���kPB��^%��èq�W�G�ӅPM+]SoT4�z�����I�6a
��x��	c6�S�f�$���:^��K\@�%�D���:�L�D�f�	w~~WV������8����/��@�r1��n#���Mk�Ѣ�h9���.�1�k=��[5B�ns�՗J]`hH=?5��R� AҬ������a����A��n_&��5.v��~b�Mi�g�*� �����>�w�"n,'�O��~IϰNq��e��U
���>s�$�	�-$�DK�"[B�F}��E�����:S�ag*e�ИEߤ����ŏ����H&�c�E'`��6��uJr�+H�C�湬��j�̲Zt��a
�� [�2���;�p-^� _�g�k����_���*v��2������=<�Y񰾮��j(]�"a�X%�+.��~�B�֜�!ӌ\Ӣ����b/e����贔��s�l�Į3k�~�zDk$��F>��b��(�9�P�&��1����V��V����	���@Km-��S�[��3|��BF^")�<�1� t]^�������m%���Q\�'UE-a^xTl����u���k�@�M�m��k$�$����-�ʤ2��^7e�$34�F[��얳,S1tҭt��*�;�9�}��*�,�mȌ��&���w�Y 5��5�"0�ƀo����=��,��k�'�Ε�&b�]u��06�xZ��\���;�2F�R���Ri�웹$�=�]ue�ev��`���ee����G.�:�#�6C����*�_���������g�ތI�`,>�E#{�TՈg��$�<��.���SD����k�	���w�m���?T)x
�eʡF"����H�N	����;Q�<��^��v�M���13̑���-�n$/�� S.��Կ�����	�z�<9e1�BT �sw���J�����>l�
$sᔁ����	^�ʉh�8�����rr�.�n����檴�ǵ�e�D��n���;�;�B7���sX4�v��>���m4��O�Ӣ�=��D3�X!$���1W�}�����Gݥ�r���&�ŋ���'k�rEŽ��F���l~�`M+5�t��7Y�TU��nC�܋ d��ǚ��@�C6����%� A�����5�����(���ŶW����K6�����RtHfW�1E����n.!�Dl��1>B��7��ٜx�f������qk����P$/�r���Swk�y�66x]��f��'R���&�E� P�6�-���{��;���Y�����N]���%8u/�yy|,'�f���X��G¤k�a!*I*�a�_�����`��l��NI��!D:@����5�#d�[����R�>��Z��Qw/z�؜�fV��Z����B�9��D�9<B��G��0�,��y�P�;��/���-Z�+!�ΘI�NJ	�GxM�N�>�A@�g��C���}͢��G��Lrfo�"�G6��2��{P�v�,}�TWxX!�{�_�����j2�H:��g��}���'��� �����Qn����1Z��eY!s�e "������k��-��0���}����/'�s��I�^����N�R����:jH���d;�JJ�������su���D�	<ع'��2<�?�A���gZ]��@�k������r&�6F*J��\� 3�;�i�s����#����=�ner����u�0d�p�L�dH9�6�i�WW)s��#YB����4�?ʌo����:Q:�Ro%��L�wv�0�B��O�;�S)]���F���x�QE^�|N򳝯������L�1�]5	C	���7iJ��E�*R�s��L�Z2b�7˴��­�N���6.�@[1P�϶�4��dn���F�sF�c�4�l^�~�3���r%m�{y=�w��z?����"�!��8V%H�n��拐�
�n����!'|(��n[��mگ�	�
a��a4Q][I
t�ͅȄn2�L�2�8W!:C�w��P=��9�K+�oI�#��<����0i��O����@���:?�t�&k�S!.�V "�*v��I��e^�(��*������}��WC����Gt&����c[ؠlN��;HK��⊣M��J �I"�曬Ɋ^Y�Df>��R"�@����v8��0�0�mF�1��j8<�[��[��[p�f�<�̴*6�i����S-��s�n�w$����̫�t`K�|]�sboX��CA�I�c�uH"p�
z�@�!'���2Y��W
����$��辊ri\*?L��=lo��'r�Ri0��������N�(i:罕3Ձ]��J������$��2#�q���}�G�` W���wu��7	:R�3J�V�8<	ݟv��B��
p������2H�V��Ʒl�2�0�j��~�2^JU-?�kF�L-ը����&��-n9���/ ���M�-P����[^��CBQ4��}�<;=��Rx�J	Wa�gfJ�=J��t���0p�����opUp[��#S�X	c������N\���AX��0�\�e�m�,����0�t���,тY3[9�GNO�W%s/�b{���w���ލK�§V�p�@�`��~O�.t����#Z4!�(�}?�Ce��Ǖ�T8��p�=_N���F���p׾��������&]G�!t���s煉���9���r1ʝe��7N���,�J����5S�I�i �3��Nb,�l�Fd"pZ�_rMg�,%�Qqo�Tp�y�4�1k�M���_E���;ϟ�x�+����y��Ұ�+������T�a:vCq����#�ո ���U�X��Y�f����0���+[z��v���(��+ob	},6�F3�Q����*�(���K��1�-�#�O5��,32�\[��tA'?
���ܟ�O� �g3�I�<��9npD��T춢����1��[�� ������_�|
������������z[ˣ��[�[�����cF^_�f�n�v��e_٧o�,��a+�92sSޓ<��*\�˕b�I:�R#qZ&�ˆ����F4[Q��?@|̜�m�}���N��B�v�-6Ϧ\�eҌ3N�}
`�B��:����]���Cߪ���u]����Y,�f Z�oX�2��_?��L�l���¾����x������.  �Uʊ��y/�RT�ݝC�Ӎ�辥Ob�Р�A�=��Q���ۇ4��I.lz�k�>�5]J70b�~�<�2��:�>�6�k$��o�B��EOp�}\`�?� g���+p�?{<.F.T���hS�=�������KԎZ�̫�0q����9�/ْ]	�Jf�pw]j�/i�8�����H�B"{�������h x,&}��}�
�e��+���
>�d}5%�P�k��YJ�����{ϸ��)���x��5�,��
���J��7X�q����s��R���)����2ҕsM0��]����9�[��`}ͽy9�M,�j�GR��)�`�1ϟr�1Q��h�"[`��/V�L���v�����܉ hJHdPF=*}.���9�!cao�UQ|l<�g{Z�5QF�څ��=� ?_�bp\R�=L;҈Y|��[�1|ߖ��U��y�桨1�5�Աc����X7���kwl.x�kŤ�z'�[`c��c�U�{����Y�|�������'�����:Bx�Xc�gcN||5L6��u �C���B䪔�D#��ø�f�^�d~�-J��#Ϙɰ3���[^��
�Y�n���D��frW��n&2�!E��6`t��aj}��Уdz�� Xۮ7;я�����\��.��Qո���Z�����4�W�m�@�
�Ga���Ѥ��\��i/�Oش�U��X�Q�����B����u��?߮�X�@V���n�q쟲��@dd���*��-��_�RW���j�a-Y�,��5�gb��y���Q��\����Ǧ�߇K�r�{�����~V�z�C��Z����|���g�#��%h�Ro�����c��`-�!jzL�V��6��K����p�CX�el�@����!rɺ�#R��O�H�7�Kbw�f�d;q.�Tv��T��b�䝆������Fi��n/H-��t>�����Zb敟@�^�e�P΄�+�6o�&yyf��2U�ZVl��=�36�Ȕ�h�;Q1~%�p�xϪ��EE�n���%�%�u�eug�do�Òo�l�0����1��d ��a� f�Jq�W� ��G� r���
8�zS�>"�l���ˁ�*#Đ:�{��a��6v������o����Y��u]�� ��(�)R��S48)P�hZ���Pܡh��n��헾���G��}�=g���39PǔI�i�E�S��x�w�˿x�5�w;�v��pKB��h��J#uE�?��bJC�F";���_��;΂!v��P���3q�$؍��T������L_������@�<Og"�E��gB� [R�.��	Ft�"6 YP�<�A;��㴞@l�k�rf�e[������2}���F�{%��Ã_�n�G-��[�����+�nnZMx���U-��}��j�!���ʊ�Py��m&�������X����+�gƳg�d=�)P����gD��_�oޠc#jK4֛�	��$޼=0o�'��}#	[��+"����-V��MM�*�`W�)��I���R���-\���q����)�����]�����xVS�`��-��!<Y��Wgk�H�Y볼8;#6��X1�����Y��O	�  .��V��j��I3����r�A��[e��8ɲBf�8�7]��$��
��{ ��C�B�h�!�9$U�N9�p���%r����g���w��~�N�a-QWC��nRzh��D��\� '�}��ψSNc�\^p]���� �1R��Ur	0]{���($.��>�j&�}!��v��L�"}�a�1���*��*� vApM��]Ay��b,&��A'X�Ւ�@ʹ��!!�@ǒ��G,[R�U=�ٓI'����Chqiq�m�(a��=���T�{��<I�V�Xr��dN�&�C�Ky�Y�{��v�w����s^$
����/��h�`�	�W���q�G-Q�6�
���l ��,�߬������#����x�_����E�#_i$���'n*���9ᩤ��uC��������1J�w�-��#9f�.��P)=Y.�1N�y*�,ȿe����z�q��U^a�,�U(>n��;@y��H:7$̓�eZ�.D%%�,eBU3�{-���*�I�3������󱢟�3�% ���̪͈��kj~SHZ6#��*��L�*Rv��g��1�$O�����0uP)T쓢�@�ԝq˅ ���-�`		dHC�G��@���,ё"�uݖ�҆zJIsss(A���K��\�5e.�������T�yf�����_}� �#tŶ��7s�	�ǟ�66�������IR9�r�ܤGv맦�>��K�}�8�`Py�4�������Yx��_�B韙
s[�f�G>$#X�^��
p8´(�u(�Ja��
�1<�E����E%M���i�� �i��+��#�Q�8�H�#"��� ��sK��~�ݼa5��A�_D�,3�ރ��CM�����R�[	<�"��_*��˿<�~S�^�7ڞtb���d�����G$@� �x�r�|�1Y�2I���'4]]u�٥ׅ�J��m@��&l��/��B�����wƵ��0ډ��٢�Qک�L�Y^�[�Ŭ���T�i��Oa�l�]�o�����p>��1|DP'G�J����ߘu�J� /�.r��V^s���C>�a�Lېd?E9��K,�JMJ��Zj@I`�����|�QL3(Rg��H�/-�>���,����E���P]b�Ҷ�u:'����I��Tk2�k�`?�UP<����&Λ"�C]le�"�s.s����1�k�(�$}�eۚgN��ք��lp!T�v�b�S�'�5^�܂@	����x��U�vZ�wȐq��w��������	����N�E���ͭ�ǆ���~�ҷv��y�1�ߦ �m��b�]� �f<�:%�0��(��!���[Tq��̘j]iz�` �}�Mq���*d�t]�Ç ߡ��D0Uq�%�UK�ɉi��#/.ۋP�a�Z=�l;
��'������j-��i������*[Rџ�������OeA����$�M�x�P}b�ؘ���tQ��&�:S�#oa�0��e1E�^�E -o*�d�i�{)^L�Ώ����5��}%���X����;�I������X�\�%rV���Z�@$u�cd�ܕj��y�<�QL�g�y�I�ɞk�)[Fa�5'�}O�;e��&���e0�h}!�n�yΠ��Y5�U��g�Ґf�o��}�ʴ#�M���*�)���ϻ���?v[r���O{�R��f�@�l� ��k��gV�ͫ+r�����	d�K�a0`�w�(�/U��c/@Ρ�U�.ܯ�~Ua
+��ٛ��z�(<����P\=�AW�^�VgT~��T��x@���}+��ƽ�8]��}L�9Q=7��"��#i�J>�wɃE��g7��`��泚#����X������ ;�᧬�<`� �"G�J�+RX+�Y�2�������B<�N��"�2
x,dK��q��W��{����ۋ�ᘘR�B��;\�7��:Y��<�+�]���!p�teS��iv&���FP��ަ�?����<�a������[�~���b�m�Pr����f
�bqъ�|{U�om��%l'�Å�GF�9�B5@����"�d�3�>F��h;
7�-�Dt�� �.�Lm�(�&[�B+�	>�d�&�U8!1z`��2#/D�<��$2����Ys[�q��HJ�W�bhZ#кL��}��[��±\�5��]��3N���P�JZ�k]�cM#���K^L{R�0_냹 ���I?$����,�D�鄱V%����1+��ClK�Mc2�j�\���a���#�����wӋ;65y2�Y�	�f�4J�U���W�r�i	��{�+'�F���ں5 ���GJf��t�o����^M�,^T�bj�g������mR�ʡ��? Xic;zSR�e��瑿k�M=�Oq_�)�Ĕ�O_I��� ��mT'ߠ���2��h�b�ق]κ���C�0F�yI�M6��Ə��Z����Pˌ��4o���ef���qϺ����I�Z��.x�n}����[�I������w��gO�F	(�ၸ{�<��ws����������}��� ���7��v�pVVI.��XP/6�l]�4��u��G���{�����]\��ӱ�r����a���X��B�,�s_�eM!����`J�hG�!�:	�����}�L���r��(�̽�����3v�]d~���Ñc��em�:�I�޸�b��&F�o���^�rW8�y���b�Rc'�;Kt������x��"���*�~�6�;\[(¥��A��N�و��U�ޒ9���L���<i؇9��	�0�H�ӕ�n0�p�8��8N�(��	&k�7�{~��A�ky�������w{�!nM�۲�P�>o�d�6��t�^�i�j(v��P�I���ޯ1��>BGzL�?p�B�Y��ϑ�+!�����9���`�gM�U��%g���6JC�-��,��Y�_ Hl�4�5���Լ5��0%C�w,�@�[�C9�!����s-Ӻg��n���O��| ����]���Ģݠ��䬮�]�:�;�,Xp�nPce��~3�����ENC�Θ�0�}����Q��4F�ΫY�K�k	&� S���f���t� H�L=g!x��"n�s�&���[�C�n�ƞf�~,��˻�� �%���:�up���DN��x���J��6�9.�i;�����	ܥ�n�#ǔ��2	��m��8�r��V8&ۼ��>�{0�a��Rf*��|'����a'�H�-���P�r����^��Ǉ����L�	��8�����f����F�Y�L�Q�!?��N��36���W2�u��%���ե�`�6���{��EŪRP�\��x�����g����T������]�x1Z�"8�-���/S�r��c���|�/}R���2*����	7���w�%��ڴ�ژ��5b�l��&��ԟ{�1X��->��D��9��f��7i#�)J�7!K��q�pM=�09C���il47O_���خϫ��E|ASCs�# �m-��\�J�H�¨T�`�A�E�K֚,�RJe�3�}9�B�2�B���m�2��:ç���]]��\��wCa��6v��_m��f���	��D��x�F�u&�-�#A�6��vM8r¢RR"��.��p�L�D�����{�e�q2���&�&�� V̔d���Z��4ڈ�E��%�[�Bd�����_���B� \�E��I\�[*�P3�%�hx�sٌ+�e;���db�p�ytAT�G��,����x4�S㛦���coA���H~�8����Åd����ڗ�v����?�a��/�h�y����j�M��<Ū9C6�Q�-1i��*g��@���	���jS�4�p���khl�c��(�%#�I��`��U�����_B�\���	�L�A}-J�b��ۓ�&K����1�N��NXD=|�k�7���:h|�Q��B'�����I�Շ�IWg%9��IP�4ǂ�i���݌�3Gh���>A�S?�i�?�$v3�g��ޭ1�Ƚ[鐤�Ύ�ܡ^�d���b� GI�R�!i��w����k<eً�e���S�&�<2��|5��v��&s��X�/�㺗��(BJ>�����O��C+XL��H�?�^B֔��щu����B%.�w��틧�&�!3,��TÍ�X���R,��X~}�EMS�*�xŖ��bfr���~S�ˁ/8�X� ����4v�|�{Oe����̝�����ՀE����.�H1X" �90B�w�S�1R�/���_�U��⇑2	��~I�5�w�561�q�2&���~s$SD)���W��X��>W��T���T�����?��OgR5<�Yd����-�ޭ2�	I��b���<�
¶��o++xV�<�q3�l�j�1���9=�"�
�*��d������C{���Cɲ�:��h~��ż�W8�[��Ԉ��s�fV`�P̟��v��O�}��Hto��ޕTV��3U+'��oa3�ڼP���j8\W=���0�'E��1a���D��3�{���I�aW�!ª4ǃ��B��&u}A�~��@��D��M��,	�#3�nk�y(Y���@'5>ڤ]N��{&^���^{�0!p�q�v��Ҝf���T��6N&�i^W������G��L���hN޴@z��(�^�9�AK�
s>�S�]A#����0�̑�N;�h�-���X��!L�-!n`F�|pȑ��(l�mP�K�;��K� ��7�$w�,^DDD������9+Vי#e\�݇V�j�\�m<�r�ŵ~ȪC@�̍pZ��{C����Lߙ�'Ve˭ Tʘ�ķ�Р5|�9i9Z���|����M<�&��S���ҺS�]}h���ȁ�U_%�^#X�H�z	98����P��A�V�r3g$̡;Wq��	E?�U~������б���;�*N	G�D�E����48�+������e�6�6Q�Tk�9D��*`�(�f�~����� 14�`"}��=s����+{��ŗ��m�����?���/���8��PWi�gx�d�K»U�8�T�oC�S��^���߲:-I����j]"XT����=O��&�q�g�,�Hً`�$@����~	Ga��xL��QE�x�|)	"� �t5�J2�Y��8+g�b=���*I#��ǥ�^M�Dǧ���{f�ȶ�������NB���E|�+?m<�G�K<��?qH���%$��'�w�6-�����A3�����\��Ԙ�|xQ�d�B7�
Rs�J8�-����1ۨ�|W�o��t��Nܨ�{��`t_�o���C	'��%�Q�ZZjZtl�6Xzp��J�j8�}$d7ٽQ˃Y��'9E"� �Vb#�3l�R�*o�غ&��
8rO��1~XB$���#9am���V�/u���X'ؓ`!F�xͧ�W�g���1m$���'r{��҅�|ֹ �������͊�&\�ö=ɔ!�����1663������?�:>>K�m��� ��KM��G��'W=�8<���ME��t��n%cGA����Y	V���r����I@xf�@��������R;�۔��ӭr� .�̗�;���r�_#�&}<���׫�>;�y)�Nb���d����Y��yu�v�_��ڈAk�1��ZX���������b�93��aq�~�U�Mdf�~���#j�)(��"(�����g�4;b�wN���ze�|�_SӐ�J�﫰�wVs�Ԏ�����~�.����-�Z:v�L��]l,�*X���9I��$�O@�r�+��`v��%ɂ�{]D���'g���V2�ut�8���a
��@��y�9�s	1�nk��b�C���M��Xv���28 ����,�t�3����_�~	�@n�������_�ܼ��
I�B��g�X+|EZą�
m(�G�d�g��)|�v��d��6&`*2����|���	Ʊ��������\�0��](�ͧ�mK�EOir�2���q��ЂP�v�����^S7r���׵v�f�GsD���iqǽ=���!�˿�q*pa���R*J��dm�L�j��L�h�;���~"�Ry�R���j�r�--���&מ���#��Վ��l+ 2��L��(�d�r=�_8�^`
�gQ�b$��ӄ��9���ӽ���9hB�}�8|�3%i�]#�ɻ5����!K���O37����c�0"�����7����t�ݒ�4�&p�HKo׭4�:.tu�5|V�K_�9���wh-�75-���{B�)�n�B�t�+�0�?g�z�'��+��ˆ�	� �)����w��Fo��Q:����s���W}H�'~0��AS��R�'e�^r%r˘nԐ?�'���VA��������'b���:�_����;�!*l�U)����ײS�4������8�߄z��;�I1���W��3Z�N�P� ��@f�b��B���C
j�:/<��v3OKz]�}�����"�Jj��:����`Q`�i>�j���ד�Nha7麺���K�5�Hk{�W'��T;}U���3�ǟ�����E^w������=��ҪQS���U9�b�/}\�2R��KL��-c�9��TѫYzm��Q�"n������	�)� 9���t�.�/��종�n��H�,,�F�Ttmٛ��y���eH�~15��*g0��T�e�^~-}��q�A_!�.\�xW:�qǏ�8d3}e���_V��T6�=w��s�1�������M�A�5U���7̧����4�1{��$oȤ�2t	 \�������-���웬"+�?,���?%�̸))����N����(i
sBHWl�p�0ʹ��Y�xҀ��?�ّMu������1��ѽǀ�T��Xs�PW���J��"�_e2;��إ�*$|(dܟ��]":E���M��Z����iuq�q��X{�B�DaKEn���O���9�t} �2!z)��}�h��$/~E��b���a�P��͍���� ~��b�>'�h���/�����oᡡ����v=��|���.�,tV ��^�F2�k^j}��k���i��e?,Ē�lY�`�56 *si^&T��}���^�6���sY�;�&):��J0d��u�����a%9Y�ɺ���;�}{7 캚��,ٴ�o7���_��uYbq������D�#t�)6�Xʳ?��|�X�a~U������h�تG7�T󩡋��9
�p���R��+	64�%�y���dЙe�ǒ$\��)Jg`G���C+����� VVVVn��պ�u�Ş�w,Mݢ/��+�)�l��,6\[���Ù�[�}"��v�pP���>d�ܰ}�ަ#?��'�pѡ�+�0���
S�	�2=��!����W�賝5�\k�o��`-ln�gm��<
d8��%sX�pm�:��v��K�]�A���{��w�j��À]��O��1�j��{�/q�]��l�SY��}��Z� ��}�dW[������v�#���䥊1�h~�V��b�B¿�s����g���F�2�G �&�<��wZt�,I"5�ˮX�!]8j����e�E��d��a�xFi��w�p4;9BH���SG�z�G9D9���_p���4e����$�#���q��Xsd���ʉ�RE�*�w�q�B&��������lf�7i���i���U�A��*�b�n�ʵJOO�W��6�w%������=J1�asc��]X&/%���$�����l<�o6�ᄙw�'���6����"�A���}���EnOz���<>-tP	�TYlx��A��]��0��1}�e_��i�9T�g����X�J�����d����,$ ��p#TKY��#{}������/I7|xj9��D�T�s��-
��^9����365]\k]rF"f����I8����px-�Q��zuf����z;7{f�]����҆mG|����I�e���q���B[8�u(��Edm�+Rz֠���{�����
ɲ؝K0�j��l���a"}r�����*�
�@Z	۸;#�5�|7ˠ�.&�G�h��Ҟ���e��\�]��/Ճ�ݗt�>]b��!P��-�M6��}/���k��9��y�/|���3~MgC=��ֻa��S�>��B6����ٌ�Ol�;���)+re�*��H�g*���?��Yq8q�ޥq���a#cy8Z~�+�yt	�	ec_��e�d�,�r�	�r�U$"��?(����,�qn͓Kae��ul&==3N��T&Ԭ�Ǉ	��c�S8(\��E�Q�����M����p.�4���LL�J�~�hސ�t[{��DM}�P�o�^^_*��� ��A�{�6�0�b��~�E��S��,�Zt��g���g�X,c�=��t(4�L�/h����qSz���3�޾n2| 5x�Pw��WTT��L�[�<;Ci}��5$ί]��"�#a��M�~Qg�,�'�r\Mg�Y;s���p5��`�Kl�v�IR�7�A�!�Hx������f�-|�U���z$��!�t[F�%����0Q�5�O�M��F�����x힧.Q��(p��h����j�{��4#��@�g��,zR�i���������ԗ�*hUP�?y�Ǵ����'r��#>~y��Cl3������LJ6i��5�º�f�wX�62!�:?����G��6��cWb�����f�|���ouuC�?�qU�&<q�y������8�HF�~�+V�Tg��ׇ�)��w3&����aT�u�j^X�TxY#��n���|Ƀ,��(~	�S%�-)/����q���%>aai��4��$�\��=�/�Qڎ�x��A@��l�{>�Am�~i���퓻�&�+�SQm��r��z��vF2���~���/�{��4�v<�hZ��R�s���?������.�	�pp4�� ����ս;[G�]����ǸwkS]�>��l-/�`9��W�3MI	Gr���
�2�K�1����Pp1�}v�x�7�V:���6��(6���{L��s�z�K�D/��T'�x�������H�o��%ĉ�%c����/D�tT@�����04r6�_yv�.w����e�@�}��Z�����0���[�|t�=s�X#Cu)�<����˒i�Vȕ�9�B�)#�{l��Y�2ޘ��|Ϲ͍1å(��t�pi�0""b���+ v�)|�;�y�|��J�o���T�웷[[��xIʶ�v��wCf��ڿ��oB�R�ŝ�h�$�"ŴlN�o��6�燒�*ú�:؜O�W��-����]���Cv���Ћkӷ��aN��P�?��4�k-<�I�H�Yo�!$$�KW[éY4v�Kxӓ����2G0�$|��@��S ~�;K��gy����d��D�ʎG�����j�[ަ���g�`A�[n�C]W��,%�M���=?�*Ma���Pm���4o]�wj,G�Cve�o�嶩-xv�o�y}87+�sm��b����C��ޭoY}�<��
�X�Z{|:_Gs��?|c���BWJ;Du�E�v*j%���W��(���֑�5q-�.6a.�_�C"2�v=ޞ�{��j�cP�O9K)�ym�C��|�K�.��{�����v���ࡿdk����41)��N=GK��*�:��{!���W�#���g���/��sB�KB� ��9�,0�f$  �7#��6i*UjSSS��"�����$��>�aJ��I��冊j\��ѱ��Bs]�_�iU￣�
�iO��T����@Nn�����Y|%EY?��,m ���0^��wtt�8��XTT�����CGq�Ud|�2a�daZ����
>>�d����� Jg�i��2�o{\�������^D�����~I�1����ߑ�Kަ@�$L�/��ϙ}~��QV����~�N�L,.&;�3��1b�񶴰�7�����g��C�5���Wҏx��urZ}:;C�I����=��*���v���o	a V;|�����燾%t^D���aS���z���R[+X�AĀ4�2F�q����VZ��)�Հ�j��Ơr.|O�e�/?�;@���lF��k{�Y�+�٫k�bz&��z+������J&u]mc�N>,py�	�8��j���12)�ًU��.����ڪҵ^������%�e��ӿ��9�?�n'��Nu����b�U�>QjdW0�����薊N����y���Tj���a���A����:�Å��zD'�4^���.�Ǧ����Zti���*�*�r7H�˷���}��l�21G1�Y�^��/�@��Òi�Z���5�M�~d�P4פD�,+?52�%:�3��vwAk��z�RX%rQ;�n`GO�8(��=bYhw�A�-���P�m)�{Hc(�5x��a5T�9���Ȓ�W�v�R�U�S=��5��lkq�ff�	��w�{���s�u���eǵ�S�g$NhR�ZR�?�\;"-�eb�1�^�X�_���ҳ�N4<��da��6���w���OR�P�����Ta�͋���ǝE����#�X�Ŭ�#^N���lľ1��z6*Ҕ����W����A+5�§���;���;��4	x��$��!X�T|?m���k6��	��N��$��ݖ�oaTd���)���Ej��Vq�bB�K��4l����(5r,�9�!�mY��xJ��wZ�t�� �]�d�2^�pB+�����F9+L�Ń���Οz��f_]UD�zU�t�i���O�m:kK4vE�g�3hNW���Y�@��@��es��D�5?�pd!���U��"��-%�P��ح�ߵZ����[IiU!`���d_��SQI�i�&qы��!3;�a��Bm	'i���"�p���l�h�W9��X^S������sMme_a���n�0H�w"�����^]����*�%��[y����Y��=B�ħ+���~H�E���f��o���z�p�N��;գ'l��PE0��$�Ov��ުt���	����z����E�}�'X2A��O��RP��D�P��_����Û��h�l��s���FޠX4.�#��d<�$gS|�0�G�O�o����������p��$����4��y��ЯV��~���nI�I�NQ?�"�!$O�h��|����dl����ѧ)B 6����d��R!*2���[������*��3��UY��ѻC6�7��:n�>"���3�H�q�k�W|�6%�GZ,z���W�#�J����ǫ���S����5�6�8Le�Jx�چ���D9إ�	H@�i��NFq��$b�Nc�-����K�^�c(p6��7��C�p�w�F��ݽ�J)��p��r���EF	4�(Ւ����ޝ�.Ь�i%ۆ��7h0d��g��|�>�p#X�����)�J���`b���Re��(�����ő:C��sv� F>�.U�NZ��`/n���ǂ���kI���A�VT�+%u�Qp���U�D&�>�䘉���K�y�F�a*7��4X�Mh��}�{]
���L����ArZ��>����;�{����d���^�������u�bD�����c����$l"[���R��;���>=�";r�/�.���K|�}����uPR��gM��/JZ<�u4��A�<"vg)�Y{P�M�[b�h[�E�8�ׯ�������P�,C�1����rƁp�,��[y��s��y%�]Pe0�p�%6��ip,���R�{�O=��ok�}�Y���6i߳v����%��F!�t$b�Cdm����-���C7La�QV`�^�7=CWc'�9��s��m�z��;L@/��d�� ���ΑZY=I��k,�3�� �d3���=�+H�g��:�Ŭ� 3�y��ǻ3�,o��<C`��ԡv��B_Ñ�Ɉw�օU��Гʈ���w>�����U�uF�n73�l
{
��8sMM�?���"r?�^	��b��wD� q�N�b��s���/&+]����B?p��2Z��ϫ!�,5���bf$���pD��7�nI�r�A-����Έ����~��Li��{���X�v��o#�*���Q�ʠE<�m�V�����,-u��y���ߏ�8�=�~ �M`S�K�[z-�;���t�pBP.`��2���RU-Z5�����c�<���	������j��Ӂ��P�vZ�e���8!�Z���*�MF6��v3v�!9dm+����h�$ܠ��%���/��	ޙ���B�'\X{��uQT��D���j�S�		��9�w��2u\��U����8��ˣ:�\�y��v��L6Y��PX>'��Y'��n������"#Ŀ�w�������qu%m��0���S�7���m�ጰ��)�*v�2�*g��H��N�N��yz�b�p[�΁��?P���>���� �͎�c�z�LƑL~zRR�h؊��+�I��.ڷVA�:�7YMp�T�����@�<����RQ���.�nFhkWT�h4r�eY�iU�D��r�t�3FlC�9�.L���̍���^�����j������ٻցVXҎ�6�\�,_r�ASp��QF��%��($�Q�Lu�����w�����T4`� ��1�DV?2~���
�l��������bw9�VE�{Qh�$��	'L��&gk.xUV�`8��e3��`,p�)��#����\%E.�o̯����Q�Q$蘊�'%���o����.m�F�x�����Z}�>��t�}�p�o�z]+�o�_���Es^�����CWoДvo�)]VU���|��(�iX9�Ep�´�G��qo�������g�5��ҁJl�/���è�4q�����B��即=��]���<j�U���<��Tt[>��x����T@r��eK3���
E�t�!m���^���2��D[�=�i{�wmo�H�:�>$����� 0E�`����:ӊ>ad3 1q���TΊ��{�>#ơ2�����s@����f�:;Fk�Glc�]���tJ1l����ҬC�6�jr.�Ծk�f�z���:�ޢd�}�O������-���38���Ξu��&�w8C�̚j٤)&�fގ��P��;a�cDh!K>��@��?�AvP��/8��>l��X�H�&�Bu���)d��,G���.	
t��\JD糲杸}]QY���xv1Sj���U.	6��޽;Y]��@�] ����͖Qhg��������L-�#��(��;d�����v̘�ŷ��1K{��w�O����ɫ�ϧgȶN���O-"$�ǯ ���0���uU������*dr%8���zU ����!�Z�:8��/�7��	�L0��?/������pF�M�-�����BI|V��c����3c�Pm�9�M*Xls���A��r�o$	�5���eP�4���}SÇά��7�=�̓X�+׎����4~�v��x~�@eݐk[����M��28��H�ol�G��@Ѓ���a2�ܙ����6Q��DH=�ͣDw��w�

�_-�Y��H����7%���oCB���j���.������%�Y���I=�)ӫ�&*���K����ܫ���	$f�z�רlv�#����
�r8�?��p�� ��lN�ܟ*��wn�P�?86U�lwM*�D�u�����T/p�o(�l�����qC��0l'�����V�*� �e��%d�[V0�=mP�e���'$":[v�-�o�C  �������/>HU����ʍ����;�|�(C��R\q�߱�������u��|�L${Kf��#�WZS�E|($J{mg�.���u�W�����mӝ|�:��	R�Zݶ��J�?ַM�X�LH=Mĝ��9�bՂ��Й��R4���͍k�O�F�m��>-|~�D��W(��y��E�$�<����	w���Ii~ϒ�+� �[X�m[W�C���  �_�"I� �t��K��o�,2ԉ�H�]���rK J�)r/��VT�V��j|��ȱ�(ʥ�J�S���1��)ԗ���&�]W�y�.��G-xb�	M���X�w��׏�?8�8>w\c����%����Q�|x���Cմ�6#Y$��WG$&ھyC�V�y��3��
�z�$�.?Z�x�KZ��ֆ��Ν�(��������D�¾Z���Ґb�/��  ��#exzq��G�ӮN��� ���%V  �P؂uHY�j\�{7A	�v��\�$�]�i��D�����P<;��|�����J�u�fi�~���2�@z�jw��q)�lB�~����h��r5_�+�+�v�f�
�s��<��^��5��	��ra7�C]W)�Nj�ű��TT�{�+��;����}�70�����qǼ ^���?6�d1�5�*�P��������e�$�ˉ({���:YF�N��l���'zZ� (���Ri����������|y��,�ͅs��]���6n�M�7��w��*9eVw�G�]��H:v��ƍB��<��UW����T�%��Z[^�~��N\���o��_X��3E���\�>m]�Qu܍TVj�`֏�LV��^
��LE�*oUW�k�� E�$�4>�`���j%Sl��>�?�a�XԷt�;�$�C9�ϗ}V���OW;"6��%��m���j�<�.P�ۈ��z9�y㩮���]2��ޅ�L�̼���ß��C0R)�w<�`ۗ_O�r�o쬿X���v�Y>�
ȋ�/��w%!��\O�Â�����f��j=b������$,������k��llIUǹv���&�4�,��D�Ta텹K��/�����=q�&������B8|~��q�#a�����+���+�F^�t'����>�jP_��q��>{��7�Q*���J��7%�ƪV/�k���~W�@NM���W}�W���3��Fd�)o�����s����9�y)+;�f��Sg�R�5�fso/~ݭsf{�WB2�ۣ�3���ˉ�|���/�z��bzCFln�¹��4d��A ]��v���+Nb��6*Z��4�,R��^c��:x��˶qzi]�@`������|��$Q�CF���e6��
�r✾M��CNi�k��峧VWiGj8V��O��7�lC��{͒����>?�k�E%Hh{�s��E��F����26m�P�7��}~b��m���(4��ĂT���7Ϩ���?�
H��{|��oN|�pL�\�7dxr��"�DW��~r�=I�
]ޫ��2)�9�כN�0�yؕ��5��S&SƋN*\B,�,o4���{s����T��3��tks9�|l����HW�.z/�鶭�m]R~ʳ�/n����������<-w^�����R�0L�֣К.pX{� ���.��\!���$2
�Kd�`n�����{�SW�������[<1����wi�@��{$�_bl������#Cm�ĠYl`_q��� �rвq�Go�x��HN���TQ�J�x�h���=[�fgd�ڧ����V�3�Q���aM�|��� $�|ˆ��A�˧0H^.V���ܡpi��T��-����K��$k��O-�9�B�PǲD;ʽxR���&�+�X�DR�,�t6�oE<�j{@��ѯ�g���������J���N�?d��S�t��oy|Sc�|�������F�b�l���"iL�Rth�*�+��2k��_����עcE��P!E9(�{�O�\�;����>C�������F�d�؂�Z̹�l"+2�֬�TN @���]��W��Y�|�lk�͡�_.�{��;O]�A�;B�>�vJko�[%�V)*۶�~�:���b<��k��z��t|c	���c68�e�M��6'���YJ;����vG�ճ��m�u��r�ut_[ ,��ƅs���
�������(4|��RM�ڨ�
�}!�?;�U�z��F+і?f�u[v����r���Qt�aM�aW>B��TZ]"%�%���ݡ�t�t�%6BJb����5�������>��ܿ�<�4�u�D��o��9}�A��2r����+{�_�p�Ó���E|�=&�:E����^) �#|��ܛ�#���$6h�N53��r��=hm||��G|%
@43��?���^�AcN=�]\° TcB�9M�� �ܔs��MV"{��=v ]��]�U����~���{�x��2<'�8��iM�r�;K4�n�4�tG԰�������>���傈M��$פ&qIo���3h��D'D9s{xG�|�cB��6��͵��$-�a��J
n�i_�lVo�^���������tN�]�Y�<�����N8e��w���UY[ -?� W�S$���O��䧋^C9��}]�Cv"�tާ�6[�%�B픥w�X�i��ԓ6�r�}:3�f�k��sN>W�kq]?���F��t/�H������v�g�}.�a�g�Sz��Wp�ǫ�:f�TM ==���ɭ]$�W�����m���[V�SV-7./����D9�Gc�g����rI�z�'��`���ٙ�#=�ﶘ�E|[�����U3j�֢_�Ņ�]�Q�<��t��N�t����*���%2���9�G���&��%�9��x��:���h��X��B�T������*b��t�����Z�o�m�(�� Y�p��l_f�cЬ";|��M�o��&+�����]���f�,X���Dg������Y�!�m�c�w�����8^�f�8@����?�*r��F_�H^�3e�
i2�I�b�=�w�������mthk1���{b}֋M�wc�|�/���Q߻Ba����sa.���ӵ�o�AԶc���{�& :��^�ݳ�� ���W(x7,x�k9�]�D7-l��o�����V� ���1b�S�����j�	 ?hGK�D9;-��f}�A�N�Q4���|��ic�0�+���P����:`-�R��8?}�0 iw�����ܾ�a���j~�-b�h�|�͗~��wT�H���p������V�yQ�`ǧ����E�-�%<��s��⛍��A�"�����yF޸_�#���G���Mx���4��Od����^�RUd������vd�Jc�qJ���yaU����a'\��`<r	�sz�~a�/���H0+px���B��G.z��u��*�:p!h^(;���;�k�:��1TL-xÁe��J�bbk7;Ԋw·0�������a�jʶo�w�5�id\�����u\�pbz2o��OE���$��;0=-��+Γ��&>�/-���-����u��Z�V$;>xR�����ٍD��-�>#�ͷ�V�xK�b����Z2�Q���Ȯ�Gа{p��,�/ErZ=uF�9����1���&���M���K��WG_�T�Mj'�{P�����[`�i��B�K"ŭ,V�t�"G7�v�@���mbF�I߽{^F�+��e�vKq�ӌ�K�Ktl�M�Q��JWO�vˮ��G+�Rc���5��]���x6���<�U�_T�1�br�@�p��)�ά.��dp$���7N����ތ��k���l��O��r����,��X���� ��Y�2kR��,k?15�߬7�9�����F�+�-�ߛ4�{��̇��J�r���I���')	7�����xH5W�8|�Y�}�ц�7�l̎4�^��q"�X�f�'�Vq���I�>�T� l�1`m�*[]aB��h���1��8��Y5�wRR��v���d~��@��ƥ�"�m�!!~Orrh�SY�9_�v����ֽ�'[R�N���Ps�W�}��f��<����Z�N�ҽ3f�����Ț��L�2�?�;�g����?q�{��>Y�<8 �>z����ޛڕh�����O/'^ި�� ]�x�!W#�_�������)����H�v����'+�h"30�8���������Zb/ǥ���F�pTF<�{X�p�xsr+}uSó���y{t0� ��^/��l�$C.�
��ѓ�5�C�'���e3E�j�� Ul&J���wx� ����͞bZ:ˏ�;�O�<M:�{�YB��>$��Z>�{!x�ә-�#�+�9bl�Q� ����Yj������tլ/1Y����	��=&�?5&u�����b���M޾��۷����1�G�J���	@�d�n$��9{t���
�v��]��Z��-����ҟ��J֑�������A`r�4X1���]@��u��: m�h5�X�r��c� �p�?
���+�h�e���e�c�V��!!�]g��Dz������6Nm^���fѩ������1�Q��������x\^M��Й�S���C\�92%bfW����c[�R�ʬ\�=BXG��a"�#��j�䈭�ǉq��_� �����$l�]�f�TU$��4?G��/.һ��uJ�
�ɲ��v�/|\���Hg��&��cA�7�ErY6Zph*}~�w�����j�&|�r�7V���W�O�i��E�U
x��/K�6�]���_�5<!�V����:�N��Fy����X4�kջ�G�/@MTLL�.Q��Gr%u�G;�<.ʚ�mϪ��PG��23\	5���������ᡨ���ɉ��p�ۦ��]"�:68�R�3�ˡ���)����e_}�_��*&{����*X�.��[j�H��
���]N�sUְ�d���¶�&>��p�2تM#��Ơ�=��j����/�	�,����wL�d�+�VmT�\�bl�~o��YJP����VZ�mkb��{X�ss��2)�33|l�����H'���oH��I��T7����I��o_�V�ȟ<jW�	�\�^Q� �uO'a!q�:���AIi߸�1O������_!צwҒ!W[>_!U78�J:�� ����\�_�����S�J��8��>Ƈ�1�7ҝ6b������oW���=T�b�9�ӗ��f�3�lx,w��=#�8M������F�P�ܷ}�;��?�Բe�.L�����R������I�Y���9�����k$J�ы��e�,_,��� �\�T�R���fg��XȲ��'����
�pS�
{j>P�˟h�׀���ᯎ*H���S�'/������<CW?P)�萱�G��O�<��ŀ2{�Tې�~�l-$�匷�z�g�Ac,~�v�Ǉ=�?�w�I�^���V�ʿ�>?O��>:z>JV�w�Q�����x~���8�x�U)2���"w>��g~������9���ϛt��ā YJ���%�@e��V��6�L���g�!Y����R���ȭ"�s�Z�Z�h�˛*��q^H����c7R�e�i��v�!/ ��gPC#�"q}��� ֋T0&�e�W��~U�U,��o�l5�uw;��T����V���i+�������ZamV�� ����7NH�@����8�j���F���c%�	}��(�#��1�%RHm �����g�u{n����J��%����mA������ڂ�
y�1����G7����g:6�|���6�]��5@���]�O38�<|۰����;]�&��1oya�"с���
��yjy��3̛Pf�W�{�����z� [X����n(Ǿr�s�w� �.9�t-���ݯ�J���k���H�����\]E���H�����ȈIZo�cP)s�$�CoX+�@������h�ʽ�{�.�	 c��T���*ξ$���By9G�9?���
��4�;R��j�Ǡ���s�{X�
)x+�������Fr5TO�ފaJ���7K-aB�4��1I%����g��{���o�?A)�D���^�����������RV=�]�S�!�!�ye|���V���b�0�]^[�ː��$o��φ���Fc&���,�.#�qx��N���<\�T�}�}Ш�ԇ�Ò��4�,�`���6[�#Vs(��O�x�]ܿ�D7
��)�a��ę�� #���o�Ὃ9���I9U�1i�I�� �(K�Y�7��[�2�J��Ͽ���lw�EgRq���/ám~��/ϡ\�\�a�dCĎ�D��Տ�O$��i1/�+�.��?�ϊ�I�&�[Ȅ��4�C����"�+����B�Ys㣁 ��g��ݳ��o�qS��a�����g1���,�T -�nͰѡ1�qT5��zf�mZZ:w��i5�`l�#r�I>*L���������SԓA$���`n��m��	  a�	a��ps�����>�=�j����C@�R��Ŗj) ���=K�~���_������}��>i���P��#��7�*뤉�]RƓ�d�_�X�r|Ͼ&�,T8�/Vr�{m�[�r?��!dLI��#k�%��vZ5}¤2LnC"i�Ù$L��wϣ#6������gk����ʘץ8�n��T�jYD���W��%ܶ��c��(ݎh]r�V3��34p��3����^���񡥣㧍+����_��do6�& F�tl�.vF�k�l��]��z��[���uLn^�{H�

��?$���H �w�>
��m���O�ச~Y�J|����g��o�Iz	���mf�?j���jU�bR�&���GB��dNj��F��m���O#6S廼�A:V�8NL�i�yA�������/�Q��t~����6���dgG������c"(�A�+��`(�<���A%��B�V#iU�s��p�6[��>�U�9�[N�^{y�3UtH����]�i�_�5?媿<�ř�ZT�M����YY(�htO�������Mܱ\w����/��s������R�'���u{~�jvv6��Z�[h��{������Q�
x�(o�������L��B��fh�P�D������;���I�O��$��Qa�p [[fS��7�_Z��׶N_����� �C�Z��<M5^��Bk#C�Z��U ���"�w����%�]�eݖ�Y�����-����*���f�2���u��d:-W7�����w����--?t!PgC�Դ�-�i��������D��SM�~��W1)�ӧOKh�,p����c�d���_�5v4��i�R���pq#�V�Ͷ6+ ��8��#Rz�Q�r��C�������v���ӕ��0O�
�`T�n�5w56�ٓ^===�����̌ѯ�xiڻR�ܔ<�lBv��s�o��Oe�p��u(g�o��Q������o���޽h��Ϳ�b�O�����g=깍�	��È^<�������?J��墓%i�B�:��$����8p��_�}�:��P�wM��QY�lˉg��kڱ'���n�7-��A��2�&���w��p���Y����i_��*RT�����gn�K�D/U��n-F�����7%���h�$�0�!�ע�J(��֖��7�q�;�"i�[���O̬�r�E��sTEe�M***�]\��`F?CAdeK�Ä�\����Þ��&^��#D�D7�w�gi�n���ի�w��u)~����Y�Qi�a7�� ��!&&b�`���£��k�Tt8�	5��� 6?u�v��3>!~p*�/�1��m�Ej�Ǿ����E�I���H�fe�S��۩|����'��^��<�j�t1��&;VTf%e��y��=��`����h������m+aP�_�c����:�H���t腺�Vb�G�w~��t��f?wH3��\�3�ШB}�to���%X��
�$l��m��m5B�U�7��R~7ǋ��N�B�F�z�@/{���/zN��@��8f��[7�;
*U�����8�����֓��.~_�l�0�X��@/ɤOb�:����L.Z
J��4�M�yd�����b�NlE�8�5��[(2��@UG,�a�vY�lӬbĵ1�>�K��a�W\b��4p�=$��oH��	'T
�/��CH[�\tƊk�y�I�K���?�3���,�5%��|wtT��L���o�"�l��I��uSղ"2����c��	K[{{�e�t�*p��}�`�=#2�N��+�����50�������X$���U^ᆕQ�0F-��1۩ae�,3t�?���)�4("x�EO8�T�B�z��_�Z�A�2����Jr^����L�jb[=éj��.�/��n+�;��:{lǁ���6R�s�ڿG*�E�Ƴ�_C�l{�\x�KטM�QUZ	�=�{K�0��1��k�v�j]�W->t�{�{lt
�yv�헓�AC�k�
tG8Y��oyK�j���8L��	���I�DL;z~p)��T;�"q@-,DB�3�[�-�3S�X��rw3�-0����o��!��LZ�hCޅR�U���Hp��p�
�^+����Ct㨲�c�n
OF[�ex�ـ}Foڛ/���p�&����~yG��R�Ƴ�͝������GG����&`z�~g_�Dv'�����G��0��4�K�Ƅ{:}N�r��wu�L�r�7��8O"=���Hmk��2�"D�F8o�Z����S�sg�盢Q\1�����ar����q��Nƞ����Q3VF\��N`�6vչv�^�d\�D�Qy!�7�I|.=>��5\�(�}��� �0��+,Y������忻���yݹ1nZe��B�
y0y�`\�N�t/�Z�K�hcgߡ]t�}Xnל�d�g=��r:�CO�O�!����ZJ]����U����X���[A��۝���k��\�r�5��1 ᙗ�!���N�?sj�p[�-j5���0��!�+GUO�ı���Q0�z��$��	�m�1����;�&;v#-i�p�N�y�~{������u�M�@tU��8�pxڂ��;9�ߝ���J�fU%$:o���k�g�̟�Ϳ5�!���L;]]5j�;��*���X:����t>��}d~��9�7���{&xZ��>'�DA�U9�Ҵ�%�nb���ȕ��Cv��r��91\u,� v�^9��G�D���'��#48�]��c_$����/]����OϚZ���>
�SǇ�}��[����iQy��?R�F�Y~�Vl74lѷ���g#�	����X���s���������p�CΧy�nOG+������YC_�%n��L:���H��+ ���5Q�`�A'�l/��m�w`�W�����`��U���C� &,q~K̉e+��a�/a���ȓXָ_�ui�/�R�/��T7�Fm23�ԡ����/?#N�T	׼N����i���'|B4���zFn�[E�O��k����kV�Az0�[Z��㮑�趠�p���m�k�*{\!Z�������%���܏�����Λ�|7_���2�>7����:���nζߪ��_�P�.��S�eX��@�Z�-ؗݡf}�<�����DO0��Ckl�\P��);7�"�Y�Fa��!U�B4"�����峃��:/���
����9�ẏ7�ky�5�s�Εc1��N�B��d�7����bP��R����Y��^�>ea����(F%Kw`�S������nT�u}��A6!U��g���40�I�O@|�.@�P���k}=���*I?^hף�TP��q��Y��k�y1��	Qi���'$�B��(küſ����˅�_�|�����2��#�{�&��YS�n��}]���F`�Lǽ�:�;b_�r��$��{�k�.Y�_|7Z����rXDs��,�jH��~����J�4�<
R��C-=As�?+�X١�vR����8��I%�����U��w��~�T4�^�z��X�S���B�ͅ�T��>����ی��S���͋�/iC%�K�oo��-~#�9_�{����_�@�H<����d"`��{�$Z��Ձ�%���^������)bX��6S�m�Ul=�3^��? �ׯ�#d�Ƿ�M]�o�m		����Y`���״gh��-~-�㌐�Z>�\[�|Ҹ��S���n��^����O���SS��F��y�O��Eb�e��]Zam�S�_�^�3�K����[�g��ZY���fv������tZŔ���CLe��ɬ���:�/��~���^��+�Ŗ�:I�x���!	����ڨՒ�K�E����=��_'�F��Nm��g���V���ެ}'������;_+�-�R	/&in6����(0}�����s�߹��a0$���d��I�Q��g�G��;��.�<�:�Be�򤂆�jS�WC�)�bv/)�p�q?mz+_fn�Gߨ��~a��D�&cZ�x2� �3|~�[hm�dEL�'���C~����B��.���K1�c����.�W[_�}�/��RY��Q���
��L�+D�0bu�|�]��{""���^�������0�����MNQ,��s�^H]��hಔ2M�a�1& 6GE�D���ʑ��x���u�.���9+[W��/������ۅ� D
����jWI�!����YZ�Pq����@���Z��5>��S�^�+Z.E;}$�}B0IVmC[L#f�|E�ܖ?�bآ�J(���)�������9�ޞ�y�X����;?��e��1�Ù�K"���=����yk���j��FP��ʲM=�H f�L��}����o�����������Q�����g�����˚?�y�����t���5�������W+����G;�F����H/��^h����C���~��#��UL"�"e���|��"`�M臗lq�ا�RH_�[[�Jz��_\��>W�~�4�[��i��/����$xLq���J,�ȁ:��2���5�]7LD0	8y;��d��w�4�����?�FX��֭��ӿ�g1+c�\�j�y��կ�&�)r��:��\n�����|�\�]�NC+���!G�a��;����+#�vc��	���h�a-��a��{�x8�*���r�dH�����w	�5�Bq'0H�j���i	+�r��1������mz��Z����}��P���,@���� �DA�fJtb0�[PP�`�χ7L���gW�����;��	�2
�CJ�y^�d���2���f��K��!���޷k��;�� ��S\��a������B�K���e�p	n�D���w������);��322�M�N2+Y@�}��pM��gg�S=c��I���ڇ����3��T�I������J��B=#�<�ȢDJ^L��� �R�=��w�s���Ȫk�k�b�5� 6N�ю�JaT%%n
J����_!�7�-��p5����X��G��D}��m��Y��*$�Hס�a#��݂��~�x}��d��x9'���7�y��������a.u4��0�{ �tpx�j؁�B���(u�_q�uB�T�}����,��d��vOk�'��L;6u�Y�w��k���9�o_���	Ȧ)`d���o�����,b��st���ql��
ǵ��|��}g�^ x��
���`�+eԻ��6)&� �+��h�ށ������8	ьk˽���,�-ө��n�P��`�AcK��i_jNA��/��WoU-�a�;gOT� �I��Sީ���jz	ߟ!'��e���ʬ�S�iXT��P����c�r��Z:�Ah����u��!�.�q�9�bjj�P�Wh����|N�i�}�d�5R.���*��W'�飊C�#�p��� �^z��,��Sx)���/��h�M(o����-�Q��r&L&�r�����mNfn/V5�[�}x�w�x4�".�e�n���2�$�z�?/���yx;�E�5���')�P�^M#4�`DO�c���NVi�`_gD�;t��g��+ M��۸�B��B��(;є�Z��<������S�
�uaNC�~ؗۄ��C2/��GY��ٻOj��"{��h�y�DH�����X����b��'����kkzu����^��57o�ů*g��/��!>Eq�d*�뉘�S�_!�������*d
̠��a�G���#Ň*1T�OU@�f��*|�y��Y�x���[��>��{���WW��e»�ć%�{Yz������Z���f�k�bQQ�4�-a�]�:���W�-�W#�9�������7��ϛLj���Nٞl���@����6i�M��@�)X&��
�b�����v���̃DD�dXui[R���Mvᡘ�t��2��z����}BX����眂6[w���w�'5��)�,q�T2U���X\�&��z�d'F�Zd_GcW頯�q!�h�iٮ�NО�x���1ϟwf�(S��Iy=S����4���+���o~K�-��]����9���a����<��G'���@��ޟ4_͠����Dg��;���E�Dܬ^i�F��(y��J_�8�/�ow��^�Ȅ���5ӕ��𞷻H��ꬨ]��8!y4�*8�z��Ӆy͍�ـ�Ag<�KL{khfx��Ɓқ,ڦޝ�b��"��Ew>��]wQ��S%�A ��1��,���#��Z1���yM�:3>z�F'� Y��V��A����h(���']�z�'�r.�Y�Ń��G�q����J쇛]!����U�����(�]k�7fj��%�Q7R�aj$4-�����_��=Q�#�,��أ�ֱ>�B�;�N�|;Ç/�~��Q47@���9�Gm��.Vd��U��;3:�/��`͠���P�����w�����ː�Ç�~���{l�@Qӿǣ����� t\=�AWTE;����9w�>��q�`�zE�>�n���m�����m &�6���G�=�����7
���_�#94f�^�ݲ�Әx�NN���Q>�3��� o�C�0)���ě��ͣ��cvN�r�.+dd��֔�U�b��|�^P���װv��%+?3�<9U�1Z��p��p,���n�<L:���o��4n�VeU���Z���8u���\O�^�U�n�FO�x��W-�݈lFȚ{�4�P+%�A�χ�S;�j1��G�Δ>I��<Pv+�mt�K{��˺���R�f=�R�"Ӻ��8()zM]��o�i�*u��Q
���0��}��4�x���j�Xr��{%E���cZ�đN����8�����`s�kBF� e1�VK>�%#j� 텀%#Z9��b����٦Q���t\���a-F�җ�;�k���V�����h\~�^Y9&��$�T^g��b�;}g��v��E�4)l��=���|*GZ�B0!�/Dh��Li�%���;=`eE�4�3��p�������EY�ϥW�z���-�J�����@`�J��׶��T�AL��J��UX�_�1�ߌ��rj����ۧ�ggo��i{���I��A���I2�r�>�gQg�{�+YWb�_��a.��[]G�k���ӹ���a^ȃ�u;�e%��&�!|����mލ��Y��]�6����n��r��� ���6�y����;��*ڳyG��������������ʬ���c*3j(i�`n�yȵJ�e=�@���L�3�>�?�*�>�%�4M֦��`:�L�zP#�Rﯗ���̝�l���X�j�&���*����*r+����Ci?��&�.Y�$Fŗ�.Cn\�v+������m�S��GfmM���울I����"��q�>���+��k��?D*qk%��:�����.6���;QU��f�P���'�w���Ƙ�ɀ�f�]E0l6�苟�)1V�cV�b��x�>]�0��:��k��TBh�+{�������N�
#�V�!��6��E�ola��m��G� ���5�f��s5�|t��x��K�{�������^J���n����(���`���嵣 pW�sӎ�#��嵺y���X��J�:�5F�VA3'���X"�9i��.ҙת��Np�kD��X;�2�q���jJ�x�9��M/xM�u��=�<�|�Q1���ۀ4�1{v����j��1�O��cBP:~��$.�~ɿy_�"rpQ�3��0�wc�q�mZ+���Mii�(U,*ey�I�����yG��s*P�:ǌa�ܢX}�2�(	CK����u+������g=|�B
T�V��/�lC��(������2���w��d��2Fd�gW�ׁ2T8?8|�?�!��q���Y�u,�Nx5���M��Y)񃯄M��m�Q���.3LF������%8�2p��&ݹs�T�z=I�Z[�=��]oJ@����+q���B�N�lgոu�u2b��Bq+��H��RO�u�u�@��|�L��2�sB2�(�Q���ӂ�C/�Q/~��k�.����ӽ��l�"�$#��!�T�.1����� �M��!{U֏!�R�������l'^ٻ������.��zi��g	Ok;������4�y�!c�z��w��M�Њ�	�"�����W�D�,�LJ�J��a2@}�V�I���-:�b�V@8�*WJ�M@�S&p��~�'�g0�M��G�� ���@%�Կ���xz���=�Jp�K ��
AԻ�i#��,���e��~��vC��}6Ϭ>ܜ�SI.�R�&�CBn^Lh�e�M	.��]��s�ONM?zg�u�`Wٞq�_tn���5��Q�y&�t�O1E4|�l�K��x��p&���:��<\tw���٘D��Lxu������x&�ð�@we�O��>�:�E��f�u@xWy�i�獗}9�R���#��ѩ͟��gf+|!N��KV���<I:�P�e������ �@9�>�������+�(Ę�z�F����Y��v��jm��P��
퀙=�|��Ǻ���vR��ÙA��/'�%�����FV�)2C뛽3�$�&}���� ��W���jY�/~2϶VФ����"�d���Tq
����������1_++^��e��^�.��y�oyu&�y����M{¬���5�;����)a��C�-""���<�TADD�;���y���E�]��$i�a�Cb����!�ߋ\�z+	��?ξ�%y~�4�A6?�>G�ݓ�,,ܘB��kXb>Ս6=��."��h�Tf�����d�2\�����΢���g%B{ܘ�y~j$t�	��_��;��0��/1R���)��"@�u��,��d�^�jGYu|⣎�J�/~�4�5=n�Rɓ�4�ZD_�Fd�>��0�+Phuo/��N�!�+n�}�z�?�yc��C7a�A�MfJ��#gg�(F������7x=�����Gd[ĸ w�x"�c�f��8C�Q/2y	�������,orԚ���[��������3z����	CA@̘o��d�`�* Ў��}͎����]�۠��^f�m�%��|Lqh���E5\|F��`��[s�jz�Sq�ӭ��O<�>���>�����R�ʦvw��Td�h���x�,�:���)Ş��z��U)�/�� >�=R�3󔎰��ZJ�j�󒕂��Z	�~d}���3�y��mZ�!OK��wy�+B(���	�o,+F���E毆v��� ��),B<���>)V�B�>���w��� B��^������9�����GZ���C�c�oDŤlZ_�O�g�-�,�[LWa�P'-8OYY���8}poJ�����ש�܈ȩ��^m:C���W
1�)I�����
�����^t���r��ؗ1E�첍/���9�?�7wR������>>�_�Z��q�Oe��g�<J�x_���e�I~SxP[3�Jwq\`*�{�;���H�8�Ξb4�G�Ⱥ�ݐ�"y��+峥�J|�F���}��>��И����n]�� �X�n��ld�����
���ͭ�H�HI��4�U��pd�l�)5٪����U����s���~I::o�u���{+�տݞ$|����gZJ/�㓤Nb~�EV��]� �� ���?�l���=l��^�D8�qW�r8ת\�?�'��NuBm�1��u��m)�Y�:/rKj�p�h�E��:�8�Ș0�5��+����xn�m���\��ׅł-�aԄf�wj�%�ۈ����t��ë�{�:��'}	R�Wka��&�dІ7c�q8s,⪊�O�t��V��ĩ�>ZdQC�VZ(�{=�6RF����m�wt�#���X8��S^���\��ș��Ϭ�1n�&?/{�9�3��4+�M4�Ԅ���N�&"%���Q�k�����)���� K���Hըx�V{�b��gQ�6UdG��t�7�n�e:5��'J��i�tBz{�j������czL��?|k_y���~@y���}k%I9Ķ���K�^��1?{�k��.��	��V�E�1˄$!�В�a�|���߷�����`�gH�Ԗ�B"�#����3�
l[>ىnv1U����i�֡�s���.�2�Bjjz� �oNxOK*�+���0�;�;�:Ѹ�+�<����0k��4+:��	�a� 6��2�b��/��{�e�|��A"�[}��6���*g��h�}��e�&�lG�l����y��
DC��h��8kF��tm:/7�t6�n�����6�������lQ�V�i]���]���=���+���_�g/���=��V�o^?�����_K?lr�e����3'����,�O2���9�9�O����V��4���[!��G7w2�+n��'�6o+^={�1��)-^��2��Pr���n�u��9���4G��S`Br�����m��o:��+��T97GbdT^�P	��M+)�J��'"��ak��Yoli������*�	�D��ƗцƚL����`��&�~���\~$�5\�`�e�j�"��e���Z���se?]�2!s� �Ev�KsN����fyi&i*C7�V���'Y� Wʭ���/����ؙ��ge[��������큳�G��Q)O'�.� <�"��]u���FE�+��)aE���b]�U?R�ȯG*��1ȩ�qe�הPY�E{2�yS���^�.Q�p4_t��5]�M��W�Z���2��O\|����������L��b.(��x�/��y?�rwT�M�h8�I,b�6��#)��p�չr��x�7z�!}�)����V����O��S����Lci�T�333�1� J ��i6�^���� e���-ͷ�����]ğX΢ASi6�:3^�T�FE��3��V��P��@X�i�
*otsm���W���`�᠉*�ץ��Z��+:��y��i�]wh��w�n� W-�#~��pQx(�mjd�����7z�����T.��j��-$�R��ۂ�$�,�}.�m�:���]eY����|� BU�|2/�p!<��]�(���?j��i����������d�i =��fF� M=��%�5�5�ӫD��'�m����{�!��t�NM�x�' ���������me%F�����3�e�����/���I�Ca�1 gv�mƧk�Ogmd�ѻ��\�����LN��ؾ�c	��A�G^��VPk���8|��&ƪT��f-��׶l�������0wy5�pI�&<0�2�Sq��������9I�4u�u��X�|Ӷ7q&�a��(dw'�eS�~_T���ӟ�a8+����D0�H�@wV�5�E���)x��� u;��T?��� 5������B7E�X�	�v��(Z�Ͳ)Ĩ� xϙT�3��2�7%`���9��2F���r�4tf}� ������Ԁx�S�uj)�8~O�=y�C�
���T���q���D������9!��b����lyȞ+_��t��'�4�����'y��z�ڣ��rJ�y��/�DN{����ߥ�g�2E7�L[Y��E�d���
=���Q�A�W愐���x�~2�*"_voJ���q�q�_;�HI㉈����@�d�E��l���W����?檱�^�K M�q�9`�����q�-財 ;<p���0y�&;9���Me���Y�K�5���)n���H�O�W�(d09��yLn�,4��H�SM�\S6�v?����bt�/���Ħ5�&��tN�Lhv�7ʠ���uN1\GJݜC90��ql�Im��2[Š���D	D/��ǄD8$7n������:���[��FC���/R��5݆%>�x��N��.�!v\O1�X� ��𤋮�S�zA��kJ��UX��5T���Z�ٰǄ���zS��8��(�B��D.���j��R,�&'�M�y��@X$��C�(�|p��{��+�0�6���]x�%8q�0��w+;� ����ݘa����]���`&}�*�
����d�X6�K�C���X�����<5ƕ0]�J����Η�Ͷ?���Sy;�rLx�O�l�2�W}�RliD`W�'W�� W���[����'6�����uz�P��֒e��R�Uwy���0����R����O�;�݁� C_�,?Xy.&sx÷cr���F��#�=gt2���i=�AK�w)O-G�� e�O����R����=��oc�I��&�.Pj�@���gjU��HI 3�#�z���=��P�z�{��~IQ�D�m�)��zB�j�E�f�Ԛ%�(����+�i�̨S.��DG�VV�M]%�W����x�?G��g�E��E�轷HtV� V��%At+���bE[e��e#z��{�����<���s�=癙s�@łц�L��{
�X_5�
a �=m!G��\�X��QaYx1��bj��6�n}QǨ ]x����0)y�R�S]��]^�3�D�����ǵgL���{�~�c`�l8c�b��x}#eQ2&�u��2���eZ$�J>�Ҧ���uje�q��4� ��p�bz��N�rE��AO{$�?kDs#W�7<�i�����բc���3��i��������+��Q��O7Y�9���b��׽ܪv�?ů��z5�j���?sk�]l���U�)����;	�}(%w���m���m�ziD�nv@��.FR^4��M6��dhG�������_��b���X_����
��o8�DD{*���^�s��D(���\v�|����6CقZ�����D4
12�`�|���J���4D���S��&oW|]�V���h���̜R����Н����vwK��ĳz�l48�C��O?M=��\�>y�E`�=m�w�.'��v���y�k%�5տ�~tʚ0�^�V�}�s�F��מg�440�*q���-��h�����+Z��Z�OrrQ�*�5��S�"&�kr���U>��K��B��5e�g����d�渜�GՖ�
Z���F}�rw��A����(��?�4���'rQG=�(�u1���Ҡ1����������=���N���z�9(�V��Ƶ�5��|s��;;�7��p%s;t�Iv������z���c���Q`H�~��,�4c�G�#���F��~R}�n�.�}TJ�d�Ə�1�g�i��-�t� ����*�gm}��]��nG��rAF���(Uڄ�W��v��K���S?�]�D����Sl�#d�J9��9g�!�f���t�f*��N���@���iHDqM�u�>;n,EB��K�G�qNT�ۿ���8�;�\���q��[rф���+t:���K/}i�55��~|ɇ��B�V�'gژ�~�����Y���3`<`��8F)��h�@�Q�����ꕎ�222�mn����o;��a�+/�LQV<� q ��4��a��N�1��C���-���� �8c�
n`��858���EB��w���KůSd��-�ZM����[�/@U��ڠQ�m,�>-5�%�EY�5'Ѹ����`�jk�OX������<9{��j���p6π�;�(�$�ť7l����)�h跏;r.�+�bV�Kn�ka[��=�ˉ�f熇/�wvD�����KG�i��iw�4�X��#�'{�&-V��޷1�(o� #eYe\r���:] �+25fܼ�IO����L�$�xkP��YKD�9Ě��S����;��[�� c�7���Tl��s@ ��#`�\�	x0�F!�r�n��`�0���h�������[-.0�<�z<"Uc�C��eh�a8��i��|�q�-^���,�@�j�5�^%|~5z�ied|�D���,��� ���x����W]@q��.�(���Ȏi�|�zy���o�~�ܹ�?��􏽾�}l�g���h��3ԝnv�rC����rC861N^F<��y�؞J44��)Q�L��dY��	I�@ ���%pWHR�����k v��2ĪOe��N���<Leac���pm��ώ^�8�0�׫��(J�=�Y~sVϤ�*r�z��C�O��J�k��;9E��LCy9�k�W(�-V3o].�E[-R����u����X4t~1���"���ڷ�|��[�=�-J��)��D�v]]�_ލp�'�v���Yc��͏ӏwĎl�ֳTa-������0�}���12�.}Sz�֕�U��8����������_�x"L\�.	�SF˖�:�>D-�r���u[��T(�k�k��;[��o4���d�ZkHX�vҕegMz���5��� Γ��L�u�x�]\+*���
4:�b�N��?H���m���R��83���*v-|� �\��b@7�^y�pz�qd�9�Z�i�� G*����ŀ�,##������z��d����}�<r���q����Zq����i\?,b [�:�.,.r|d��Js�RF��"E�i}����������1��wK�KIFy@�K�7y��s�ɢ��>�z��$�֜�SB��"e����#�.�J����dE�Uy�Z��Ï]E���ZZ9v*x����n���y����ه���x��C�F����	�k8@�&�+ݒk]g���Y0&�*Ϫ���oi�A?��>���o>E
/���w�l��<,��w`��C��Z-�(��i0��S�]ߔ���Z��s�
��G�
u��%Z��R�o����WN)�Y��L�k�^#��AA]������r�O��{�;v
����IQr�7�$�kʊ��%�����*�����+e !iI�o2���S����L�KP{���g��7�'��ksށ�����,N��@�S��?X���G'��Q�w���[�)ZR�UQ#k0��ٙ�5N���f���i�J��^�;��s�.�F$r���0"������eݽ������ �-N4�!�	�M����X)*,��[xE�h���šh�puR0iD��,�Z���J�m�06����E߲�G�`�}n.u@��"������u��u,�}�S=8�̄}`�D�e',���sL{/�T��[���j�?�yG�C��>u��cF���`)�6�{��]0/�Dկ�@���mp.Iߴ"}d0%��\ ˞�2.�rU|CEA�Mb�U�i%����}��oǡhc����x����8�IU�)�� X��:.Ō���R�x��D�o�o��i���T�F�M+5O`2CB/W���9�Q�䛞�<�~����$w��6���M;q=�nPR�5��څ��)Y�+�G8W�B7�������0	f�s�P p^c&�����F��1��}6iھx�� �~�§�o�ȋp�����l)'^�F�����^�^��"���_{:W�ojj���r�ߞ6��zʊ�K��Ajjc�M!�\��
s�)i�9��K�R��+��>�(%L�4UG� �$ɔ��|jӮ[V���Y�],��3y펬ب���1�}N �*Sϱ�m9y��)�Ik�5H��c�wt��A��gx
��<n
:k��|�)�6�N~|R���N��Q�*3난(���+���4n�U1�~�X�������3	{~�D����ևz��ntD��4{�W8�f��f����,e�w`��k�ku��@����~��R��v����^N��$��J�������0/�$E��g5b��康��bY"��"��͡�9�T��sk77�@�d('�Ԧ��(��?�__�Mک���Lx����ʊ��Y��;�f*1yY����(4��}��ނ�{�77���o��h�7��{h�F=�+����G(���"�)�OK1�m�B�(�X�`�}��<�/qpv�p�P��S�E��/촉!8��k2�y1�ƽ�ju�\���R��r�>���A����)�wo���ie8�G^�mOդI��H�2$�li��e�f&�T�},�rh�I:;�W3V/t0�_��ӛ 6q�L��C� ���c��U�O%�tq��ε���p'�Ӊ�O�󶎳l����٧5��_�E6��$Gm�a�1;%F�,�2�I�����?�hʭ�:���7�#����X��b� �+���`L�<f-(���\��ŊV�8g�KxU�$��"!K+���P�N�3�Ցn����W*�^.�c�OGT��;����� �x�x_�N�PP�㟞�wܜ�J�����7�^�XB���T��:y��u���hG�W�ϡ���͸��T���/O�4��@v5@$ urZ�t��4;1Gz��3�_�U�wc��z�������XV�C�W�+`��?�I3S����=���k��\���3��<�EH:V!�L�6,K6�޺-��җ<zbb�w���{�i��3~�n�E�>�}��O�M�=��c�i�0�?�j!bңܑb��uäO���Jb{��js����^��=2���	)�Bno�xAN���MmM]є������Wn�N��7v*��Qp�Ø'#��6���rO>wK4�4�{��]u��a׮�V�IYeee_���6+�<#��O�m��^�L�#[��H��$��j�k�����Jo�5�l����=����	�Ei��[ӌͿ���2���~�~����fz�q��whV��Z{O��]�+?��/�X��ۻ����'Xq�"F�Np���n�C>�[v{���]���T8b�C��#�o-�5��X��rW0�����£~\�n����/0��i���{�W��m?:��0�O���S��<e9�xS�y�(虏��j['矴su�/�*>l7H��8Kp0�rq*_��� tr>nl��2�ތ�e%����9ѽ�w�4�ªpp+�ąC�M�ᙻ�D���Sn�}��h�Y2�(�m�d]��G�j�>�N�A��[w��X�:PY�ߡ��&TD� �3�矗_pTҜz:�e-N�ƾ}��W�P݀���歡B�"�!��a�U�g�'v��ՠn=��z !"S���q&��9�	�ʃ:F#�I�� �J�Q�nC�vo��ٳ��?����3�ߠ��C_���@�g�����dJ������� ��W��a�杭IE1�HF�Sӄ��_ذ�QW����{_��"�oo����&�����5�����/�]�.,L]��@�/F�R`�"�7��/���T��:ah<��7oR��4�*�1G�!&(:ӌ�	���d���Jl������Y��W(j��jf�!�h�r��x�OX�����lZ^��L!>m]N �-���1=���O���c	B

�-��8�7b&��ȇ:�~��ZU\Z�"-o^�{~A��rT���`.ޭ7�L�WX:[�����D���ǚ��(7���NN`���o�꾾J\�āf��*(,F�^}��H�tr�f���i~=��30����.���Iv̉���ÞRF1�3�i_A��~�{ן�����(?��ٻ�6�zj�-�Õ��ry�\�8���~m��MmmHc[
��ϣ����x&�����,����b'������`�}U��B�a"��l�9���=|`ln�r*������p#���'6x��D��k��<�E\+�D8֖�������A�F�P������IKQ�����G����AA5��lK ����&J�3U�C� '��E%F���&���I���U'(���?�p����V��7�5e������@� ����L��0j�h�~Y�O��s�y���ܞ��x���O�{��Lr��B�������e$�	�?,|�����8�I 5Y���^Z�R��Ny�?
b������o��.���D,|s�"�����)���E��4f�%A ������;�S�+W��}��CH�l���WF�J�����ݔ��ד���l�䜤�*�~b����)ֻ��Y�"m��ܵ*lN�{]��er{^���H�%���N�_��0�:[/N�Ki��V��a꘧�/�,@�'V~�r����,� �}��+��jI?ҧ�+�H�2��n\������CZ?e�����ۑ�q�������P��v��}�=�;�5�^E�~��p!|�nm�����Gw�ʿ�v6 /�+�u����VX?�q<t���(�9�7������˶$�+�I�M���W1-���}�4d�2&�s���{Ҷ�|���=p�0ꢭ���u�P����$�e�wL;o��y�����;=!��9��k� {i�������6����ġiy�*�v��s��a%"��34��o���wĽ���l�ށO�RN+Lh����!������薠ۼQ�n%$b�5�ɗ���O�
�̞ĤY!����#P�2�W
����w�{ܬ�h�[�C���Hh�6�d\���P��R�"ز��C$>I1P[K�ƈD��R:	g�
��ch����&�����+
�~1��Lķ�ӠF��w�2�Ĳ���u���)Ρ�(TW�ߣ��13�?�6LV({���7�ރc	C��:Z�h�m�)H�sC���հ����~T�M��+�/���zA>��^�w$6����?� G]6��lA�j�Ku���ĉp���:�U�n�E��p�q< Z � $7��g�JE�[V'�&-��?��~`����Y]�3�TDGn��}�� ���՚jr�J%�.<r7���q�H�(�l���L89@��<"�0~]��k�|�d5��ȑ������L��8ƥ��d��:� 
g<�<���$�����g���zq	��Rw������2l֪��H��::X<ͮ�6R�WN)Y����ו���� �h�cv�� *Z�[3��9�x3vL	|�;�Ց�$}.�f�N�}8b��1����K�G�3\>��͢t�Wףbw5\m���>�!���\T��%5�k��w|��¥�o���eZg���e����'�j8����[)O��3���ٶ�j=4v��٦���!�]�y2W�Xۄ̷_���b�c&i}+�&c{/�h�F��ĥ���;Κ����;���9���*,�v�rD� �Yܲ�m:�Z~�·��n�6���c\���UVdז)�i�uG3�b�?c�w��Ԡ����O�YA��q6�,�s�`���������o#N�[�)��fD�U�$*�[ſ
�
Ԍ�X$P��wU�K�!,��^̡ڢ��0Z�Y�b!�,{c ��o�.�p �ډ�ǚDt����/"�U��Jߔ��#�f�9�����={�l�}�cZ Ļ0��F4O� �!Z)N#�n,u�Y[������r�@V�^W+�++=>X�*�QR��d����m�@�a�
.!����BHAI���̹��s0�W�H�Ɩ�d���Q�G��i�v�I�P�V�~J&�80��l兔v�	i��і�����������NB��4�=#MT��񺭶�B����ץ���m}b��PqL�~�:=�o�3S�dӦjdŴ:sN)�y�H����.Y�M\�����*h3`Y�C�y�m����]Lz��/'�'��qtZ���H�(�x��FJ����$����k��5�졬;��g+��\�6������i�A���H��8���Uy���M�x�+��qC��o�t{�����ę>�� 鍠,�3[�^H�x�@gЈyNF%>�ţf�ߛc��Rc�^ONi��
맔�)J��걤öZ�����J��#�Co���}���#4���������+����@�)t����@lB9���)���N�b T(�˲H�f���N�x	�$Kgf�E#TdUa6��B���3�����˜�3o� �%#�u+��@o~$�b�6U����~֜�-�h.
(RM�]�|�h~��Y=&�b�l�@Δ�� `(���~Y7dLRVw��
2I/z�O��o_�N)! �$��?<03�� @������a���XPD�R��'n��hw@bI4��W�+��|Z��ܔ��he5�z+5����Χ�x��N:�e�K-j��x?���.�e��2��0B�JU��?ϑ�ilj2vln���oMfH��ه�FF��ϭ\h�P(ܶ�������
�\Xx�O{�����KT$J�B�IY��pk�s�k��O{4<,*��q�q�Im�G|�G���󰾗���Do�F�+3��Ko����n�]��PZ���l5��Y}7�K�E�c�L𝳭l�>+��>��iݦh�)(��I�M�M�_�çQ*���Զ6�/���8V$��}�_��ˍ{�ł+�)�A0�O��	�L��HH���a���v��"���pж���'8@�
�,�&M4�dM#�;F0ǆ�4��i��,�� &�S{��K������@͞vD��BSjjXeH�ztո��D%�}PP�B���U���^ƥu�6HE�D�/l�6�6���\XAe���K��N�w��������>��s�]�fv	j��񍦵�ˤ[O.�|�Lyý)b϶�(�A��C_��q
w/�e��
H�gz�n3����&'���%��nZD�Rd{��#�1Tx��J��$L׬����c;�� ���9��X@%�M�/����x�,�� ɝt�z�w��
�-5���>�]�������S̈́�B>)F�B������E{X���c�T�q)� O^�K�C&A]�c�����'#d���-KR�����OU�Y���h>6Z�����з����ː�3%���q�Ζ���"����ُ���J)
��~Y�!� 2�:���O����n����oD��̎��4{��RA}��O���}��mMq�)�R�چ-�s���'�<�C���ܶ���P��[���o���Z6"��z��g������w�6}�.�b�Q?�o �N�����n�pS�"k���hR\j�C �u�و���N�J��y�}�s�>����N��?E��r�\lO`P���E�����n+}<�ؘ��ca����`a��z�6)�ch���~ō��a�N��>`��@��Q@��p�R���E�G�dmö�,U��効�o�v��a?;:�**����5��}O
'F� ���&$RMF��x�4�UFW1�����`��:��\��4���eȐ��A,lnjn�Fu\_+��i	?�`��I]�s�><ϩIђ#���n6:&e�=�S볞�^��+��s�#555��p�.*��'sFŖBS�
��/7��i��s����`�߼��K�G�6�ci�����%�o�t�FJ9K�ن�?�j���mVi��#��<�SL��p?��iz�k#։��۶3�G�m����h�XaLNp5Bʍ���[B���� �͓���'��痗�ɟ ������g��u�:|9yy� �OL3Pl@IP++��ϫ��Y�M��wZ��n��x}d����t��Cq�a��{����=R��T��x{����Q��ηr��:��+��4O��Bi ���8]�U������xKfص?P����7''��ۛ3n*�_�- mx��`7.Ȼ����K)���F#�J|LU��9(E�)�[�n��V����U��a�垻����Nl��vZ�g��>��c~Քڐ���_x��'~%%>���ˮ[c!|�{�� \�/��(�13�p"�?���	�q�>˞��j�}�*h����hm����[vM]���j%ei)�Fxz��_�\'�=+/�r{��'�mH\�F�)�K��1	�e��$n�_��=֛uzZk�^����ֵ���", t[Iq������>�	#��fEU��g�{�Nk�ƶ�N���:�->�(��0�ڂ	6(�� �A�Ƹ�E0#c��'ڸ}�����ΧO~����Z��;W��1��XK��r�å��2���\Hθ����4��4�W��V}�/Zmt�T�����Y��0�}5�����ƒ����0���F~'����Dw�����G�.��ƀ)�{�)�׹a���\��|1����ద��d�*��\-^u<��c~�F���#)J���@�ͱ�H�����L��6�4�:����fx���<kl,8W��2lR,������N��6�>�(�N�����k}�� �%�G��%Y1��MX/X�����f���W�Hn��V�3ϸ�q��7H� PH��i;F��Q�f3����鶯�j�o�o��4#g�~6×�9lD3��{o({*d��k���kYXsA^����>V��i?[$�9}�H/����ں:I���nI�?S;3�K�L(M�˪�\P.����T�s�Z����F0���]C�����W�n����8��n��������<G�$U.�\4��8;�݇APc�������s�VX?io��%���zBB�:�W����O�$L�c�I�揷��k����ԉ�Sf�u�2�����H@߿������F��3�Z�Z��)w��q]��cu�)�;����76�-�d7܍VGWw��i|�����i�^W��\���7��8�%���/���	���؈9�[P�Q�_���Eu8��3�$q'��9s)������}J�/��I�>������fjh��]��wJHS����� G� Q�k��XJ�͟�<��dZ���ȱ3��2z9@�E9���i�!F�ͥ.V���ݛ��<*%�ى�}�Ms/w�<(*`��2���E��K�}ت����&�d-�b��j��9=�V��[��J}��̖Ͷ!l+i.ؘ��`y0�p�*62�0���\f�l�v���4��B"-�%��W�52�a, / 5�G��d�~�P�0���������?X��y�i	���;tɢ�t�r���gb�pt"2_��RB��<�䋙B6��G��tt��h����h��0x�o��r���ݦ5���C��ex@̬J"�.Csk��D��}Go��^���+���(-�@8c�4_�v�8�Ca����k�~	d������q��c�!
6���b���d�=5ޗ�_��H�ėZ=| ]�VR+�O�U���8J.lw�v8�MM�n��L[��v���X��*���?L\;g�*Go	y��\��8hD�j~y��<ϫ�e0Q��Q�-�'yzW�Ҝ2R9S6�u�iI�$X?�14x���:�ΩoX���#WbA������c)�+��m �Yhm��a���T��H}�寵��w���Q�j3�F$��W���uR����agD�$��<�0:�,p����c]�%����]�1�ZP�
��.C�?j.I M�w�e�

�
����y�.喝UH�OW�.�:~4v�.7�sw����B��Xj1E�AL+x����Ͻ��0��8>���Jll�>1�\�/�O�6m�E��ؑ;ǩ1�_�Vj�+�N�侕'�a�<���oX����T�2�;_[����:Κ�N@b,��8R7�x�d]��k��a@��]�lh���X�����)a�C������\����#�AUgyˈ���)S+�CI'�I�Oڎ�l�_�9q&
����;K��Z��#<<��K���5�%�iv*� �>��?��jT���/[����BT�*��@���4ҝ̹�~5���KAL]��F{Ɣ���FH����9�3z{7%��n��j*4|�ӥ��Mҙ�P*��a�����v/����V`O5<;���D{=|3�|I�fQL��4�&�v�͜^�u����Y��M*D������w�-���9�o'U��L�7��3��2W'!Y��Z�-��I :^�a��,���
�*�b�"^A$.\R����>�UN6�`�+T.�K�;��k���G���.���OE=%R1{f��lZ�4�}H��y�no�e��I�wډ����� /�
��o��JKiU:Z��^C �Y@�ղ�m�ǂC�MX�M��O������qc=���70�UYNh�@������^�;JƵ�ٓ<�~Ʉ��j�����.��ѓ="K�Ôia�U!kq�^���� ��v,�����j	i��x�2
wZeM�Ϲl���y�.� ����O;��}�yߑ��C]�ck�OG7_ais��ps���$x?:�Z�УU�ONҵ9��b_�cx���֨� k�\��������ߘʛ;O�$%�I�����8Ծ6�2����F�F���}L�{�i�)0Zz�V1Q��X��3�'��v�+Ո~~E���;|���X��]=�Y*�^�]�����������bR�;�o�͸�������>�j&̿�oI"��4����Z�@}�q}���;����Q��ǌ����xa�q�"e�v/�����&��WJO<�n�S`Lͬ�]|zjd�QϪ�tb�i���F��B��r|���u�9�OY����{�v_8먫�ՠ<w�֤�nk��/D��߮��B��&�O˸�(PM��F�t�~���C������FN*T�nO-�J�Ǔ&��C8�80�Hj���wps$���� ��e����>�Ӑ� q%?����Q���m.LO�I�qt�G�m����֦k�0���ZT���o���G��!Ov}����B1 :�O�
ڻ���9��)	�����?8"�c�-�6�/3������#)�J�2a=OgGq�h}�>�%��vǞ�Ei�&�E��{ˇ���4rk��=�*��8 �k�=���]l�����EP4������_�b}$!K
�~�a�׭G%)T�V�z�$��@K����˪���ŰD�R�e�	>��sq�FX?/��V<?{-e] rmcK&M�>�y��{�0�f�`�,���˗���>_q�m�SHr�QcSp�����V�Gy��8U�S��=�\[�_�P��I;[k��.W��N!���u����De8��F�G�Nx�5��j�m�q�2J��D�h`����a<�����Ԣܵ���5?\Sx��eуRF8;ُ�����+������q��4�sȀ�0��A���E�{o/7�6������C�]�8k�m�wR�[y��l����I��:̿���Ma(ф�~��	eL򲶗����#�s2��׷��lF��LmQ���&�3(�/	����s�H����(��ט��'�K����^f�y����-���.���S��g���O�J��q���� �M��-0����M��	��z] �)I�Z�1k� ���ù8Y'����S��R+̩�Q���%b{Ƃ-��2cL�-?�G�Ӑ�q@^�k-�Yx��x&Kp �/O��mM�[cK�2Z
�9VIG����G\�ž*A�<����U�D3�f����<�c�~{�:�#m����g��p�{l'+�Ѧ�< v��h=d�����kK�g��1�=�P ��sH.��|�W��W�ܪ'��q9|�<�)�:����{���L#�'\ ՠ����i	�mｿ��j�����.(��� ���gF'�J���X9̍KhGտ����ݑ�>Q�������>6^�Q^}���ƹ�x�O�۔��?j�����m{����t��CU{5��DU0��oʢKܓE��>�t3��[y��u{�{��7�H�����u��dT=������%W"6@'d�#�e=MEc>z�8���(��tp�Bzq���c��GM�d~�N��r���p��KRDGG���z�Լ��/yͺv�N<^��{�*æp����zrE%o�v�����q�k=��V֐o���8b��d֊�li�kC��Y�_
-
����9����yI^q�T�}�:�n�����6
u��@���y���>��J?���Y��<~#�T�ʎ1nƫբ�
>��:C�_Me�	�mՔǃU��H��w�8t��yd���f���
����5�@tB�$��<G!�/��8�{G]Գz;�"�b��oaJ)�����N��1c���zv_D�S���OJO��;�rp{vM\1ISY�P��TH1���rxX��$����>�iU�b�|�Y�P���dM��4#�7����:�����k����n�M��/zfV}Z�����hW���;E�Ŋ��'j}��?��b��IGˬ�S����y��
���K��p}�#I#`|����F����R���id�.�u�<>�G�Z�Gy9����U^fw�R�fע4.�3���1q��p�/M�3��2ÇA�-�7�Fi�S>>�eޒ�yvY��Of�!�������`卝Ѯ�@M�@e�Et��a���h$y�4���(���Ӷ����^�]�u�xq�%��vMH����Ǚ{���aS)k�\��<�:�Y"r�2�9�Y߸�[`��];�{jWV^��@�@*v2�e����'���D�*��]�&�ͅ�ZP���}}��92C,_߄���� �����z��v��;��$�,_u��N�����dcٿYv"����?,��:m�>�eѷ�ٖ����	���)��օG�$Q��6�����oB��$NT���G"��I�`�T����J�&(��T��B(�4|�}̉0$�N�}h�Q)ke�T�i��mbus5*��J},m�u�����B
��BT�7����K�Q[����6�G��8������xӫ����pnȷlz�;w���W�LK��y��S9*΄߮.�f��m�'j�1˹}� ��T�X�`�w6d�E����^�%�-��lJ�|�l���9�r��B0��f��j������ �.�8FM�u�ěNwZ�K4�.��Q{-n�\�筅�G�I˫K��[�!b����[F��v�\���/�}R�	#�R� �ڙ}��!g��\��4��!�:ұt@slm�x�����n��b5��% ¤rc~vJ��Q3,�Z%��H�< *p���H��4�r/a2^1bR!��ڝUF-��2��I��@��������Jc����K�]�0�Zi���Ǧy���Yފ3z�~��<��14;�G��u�����E^�JMy��g�P�Y�Xm�[g�.HX�����0����"Q�~}�L��D悯�)��
E����F�g� ���p��D#��H���H�V��F��\R�]�_*�Hˏ7�ǁ]���n��~�4�p�\��I�����t*�g�vu�׷�U���6̈́��7�Qh۰!م�+���ɪ�p�Gז�y
���n6�-��O�
��z<��
?�$虜�g�{-c�	`���� Xp�dit���z;����@��g؆N��̆^
$�xޛ�"����YYYl1-��,;��&���tc>����R��k��>2y/^�͕��,Ƌ��>?�Ч��{��"������v�
NN�������?�������Q\��OUV���&tl�gb6�]0��[$V2X�,��V�0|��i{{�&#x���2�\��hL�q���=��[d���a/0O�W����fE�H��u&���q����έ�ϯ8�)��-�? #��āON.Y ���߇���\
�K:���?���S!�aj�r:{I��q�����K�z�������mߠ;ʝ+ނu��&F�C���U6�#R������̡���q��O�Oegmm=�9e	=�[�܌'s<�����"W��1}0�~�5�Q��bx��HDK�R���n1�߭=?#�}�ۊ�@�Q��R�>�w����+�W;��h�{<�%.�d�`!��F��$q�F��ݰ[B�-�q�a�񴮅����CIߵ_?��yY��lq:)"����_x�DEE��V�l�t��4�zzК���E����[/�����#�[���@k]�gZn��І>/��Z׋�A��Ü�_|?�%�Ucݦw���@_���fX �g{�w�\bF���I��患"]�\��;�}�*�Pe꟒l�����{��[_�n{/˥%xx���d�x��|�l=���u�I�乼��pX�!΍�>�W�:	g�1����?�B�:�O�)��?Z�;��V�Q�5������I���Y��k�������rh��j��.3�
��q��6]�|�V��<�Aw]�)ک{2qP �M����|�%�c���A�nPK[���Ƹ��f��})c�;Yx>M�f��"��?��C!7�E�c�<�
%t�����r��P��ͽ�Ε"��]�� �Ԑ�iOS�r9����;8�!-a���J)�ր9�y�L��B���%^\\�k��Y�|6/o�Ad�!.u����y�E7��'�W1qF�iNN�B#���{��˸�Nq��G������J�z&�K=�R(3ae����2NϦ���$�k~��X#ǀ�`QGd�i����4#�㒭E-�����_��)��g`��9��Z��	���+�������2d�����}m�R
XZ�hp0��O�
�,=&�(��N�/7����'���	� eӪܛ��A[�� �4\Z*���g�(w�/���M��4�%@7nU��|#}�t��n��4�����?C���B3 B�D<v=2�����%ec�q���~?�;�����cfT�-}r�{�K����,R��$��__���<N���i��n�ШD�tz79=�/����?�5�G��s��l�D�S;��M����d�1�s��	���Ml��R��"�����+L��̾s8�������w?���B Y�u��-�V�y	@�hm��,#M��p��R�׌/Q[(�����ތ��p����7����G�s;��}x�aq�}�$t�#�w,��� Jj���*V�N��z��S���t�����ɖ�ۺ�Q�Ҳ�y!ߓ��)l�̶��ś*��_��CMN�e�����_
�]@3Y�(b\s0;/�Fb&�$�����Eh�o��VO��a�w�]�܂��Y��6e`nG� ���YW���V	o`rKS)�#9�sz��~z7���Z��J�TY��Qps�Gg����q��	����N���]�C鐐0:% !�aRN8ztw�����|��9�:��>�}�\���\��=ˑV�o�|��X�NM�N�B��e�Ç�p�-^��]��1o�7a-��V]��*S��e��i��:sA��0��޸\���^�Y-�4�;�t��f��'7�^�|Y_"�̂�ӟ�!E˭�@r���O�)OpUP��I'�T��l�dd;��N�	G�H/՝���Ż�a���$�+Z[���]�噢��8�K���uM�����l�"^Hr���O�����ŷ[�"/��-/���^)-�n�R79n�tt�ߝt�g���j�A|�%���f��Դ5S�HR���kQ
LD�re�y_1����3�v趒�|�D3o:/���z���:K�s������Z�/���lsĊ ����Y���M.䃝)��DC�`�P���s.#@��73���k;��x��Ǡh���Yz�����ৱSʗXܭ�W:�ix�g�<OA��}4C&С���^��oPg���Ё;Ԙ�1e���ڇ�5"֞��ɔ
Wx=�g��w�ʼ;�/��-��p�PYo	�V���SDN�Ϻ���LĎ:���ju�7�a*�{!m��Pf-�7��Sy�}�<�����Y�n:��m��!(�[�8��I�u+���1k㸭��~�-�p��#��R�y6��r�my�ҶH�C��R/i�����1��اg�S�����������B/l�d�����8s�ň�Ѓ5��k"�Կ�@�@�յ���qm�/L�/R�qrs���)����]�m]}߼�Č�
	�_G�-_C��}�.����2"��_\��~�Ҟ���PB����������3�.������li��^�a��T pG�NM�\fp�I�ȧ�O��N�R?��1>N�j ��7�r�oKE�*�:ѣ�7b����lf��)�,�*5���v��f/�fH��?��c��
D�%�����,��J���籆t=a���#T���_�-\pJ����i����]�֐�O�j���QT4)*�г���{ �+&����U+2=����8��wر���w-�v�Q�����T�m�����H�M2�O�M.�����.9;��Ο�ǳ@0*�op�z����l�6qB��v'GH�� 5|�ŗ ��������D�^���6���Xz6�#�'w-�2��o��j=O��"����N��k�r�݇_?�k�����'�E��$ݮ��A
~���9���Q]���7+g�}�B߶Gr̾sd�f`�)�`O�e�?\��>{�HRQ�W �dK��WM
dpxTXߍ����{R2f�2�I�P��L�*�F�ǩ�T�o�/���C㮍ξf�II-f�zX,�^�p�y��C;h�������S�G*HJIN^^��ۀ,��흶��"Ld�D�lX��c�}�΢��M{a�c�oϖ�O�<�
�>:36x:+%ع�'�)���!dA�jх��ϙL��9���:���D��L�zֱ'�#d�c?�Q�S܍CmԿ��޳�Â#mp��1�3�����al�o+:�=��ۣ�-�A�4cT��B�h5�;�)�A�R,h[�̭i�n?<ak%>��/�[ZZҜ����, �%�CC���,��g�U>zzzF �A�*�VR��%4P�B�X�շ�t�^����w��cx�����;ba�܍��x�E>�M��eP�����9��!܏�&P�����"��>=�]&�V?�����`�BH0�..4��[��N��z�/��]�tiNLd��ZR���$�.ç7/�[�R����kB�b(	�L�]|�2����V�	���"�qqut��̞��Gl���� h�ow�-�p�<��l���j���b���<b���J��UO9��jEz:���������-����#T�A�R��)��E����X�f�0�Z��\��.jl��
%]k�V����UD�qy�ڟ���JY{,##�	-����R?��w�o?spix&�|���Ak��`.�>�`���rKc��fbH�5M�-�'������Gg��t:t�{C�l�R��ڴ�o�j\��q�ŌRGI��%�[H	~7fʵ��V��ԖO�UY{��vS����k���o����q�&g�lYU̾L��rfzr�rd�{���j��s76�o�H�Ib�|����ˋ_��L����������Xq�|�o][�b��1�u4d+�4�Ƣ�Oؠ�WgI�OT�/۪+RG]��C��W宇U��/���?������N�!3l'���̓VT�,�A�;�A5_]2���k� Bw"w�Uy��Ïg�Ӧ5B��|���G��ڷ����j��$.I�mr�L�]�GnR ]w�1?��T��C�Z�{�hV�����h�V��R��G�2����pUNC�;�t�N̡=ʧ�  (y_�9j�ޅ�<@�KZ��{5�������g?���
��)C���u���e�z��eg�R��J~��L�D���O�a��~NN\�r��rr��!^Z���l&xz���l3���$>$����c6}�\���$�up#���C�X(3�1Zvګ�����ݱU2r�ǻJ4_bb���ܽ�6���8�:B�f�\;$nׄ�~�����������)z,�?������߷
S��pg�qb%�sr�S8�"�ܕ��:��}�2���(��$����ځ��h{�W�דK�K�7}�.�������_��Be�y\_��ɜG�u�2�ydj#	ֈ'���ڇw�YinĖW�ES�@ʇ{7SBO����XB�w�Ts�MoY�]����뛓���2Z��T��,�%Ŗ�m�֖�Z����^��o��g~A�>���[#�1�ʻ��s���+��ϵ�wm���I�� �u����'B�p���P��}�Ԭڷ��Ź�d9�nc����a��7{Z�-3Ҥ��]c$�)mW�����dM��F�j}L�V_�}89��Z��m�g3��~?�&rş?��g���J��̏��8�}Y�y��>�׾��L����<��v/)3�p�$P��,��3zS�k�7��I^�' 6������W�o��n�?�C�}%���<痉����@��_%Ǖ`x�]���S�7G:����fzj�#4�[�Ԡ���m
�to1M#�[i\cڈ]�z�n������?�b�O�+���� 3&��Q�+d��F�&��h�ۤ�����/�2�t3��^��E�q���\4�'��,����=q��]3���_����	�tJ���d�K�5n�v�w����쿚�2S��t,�_���w��]l�:�G��c�0�S?�U����Loj�?�%��JjX�A1��?�3,���;�%w�`�b��LG���|�N*�s��?����W_�A-"��><��rT�'��'�z/ø���	Hx'��J3�
��9��kpQ�&���`(��f�kݙ�st��ݺ.�p�ǒ2��WV�P�Y�KA�c؜���|4�o�A�_�,P*W�f"u%�KM�����b[Xur�}�̭}�8�嗞YǼg�	Q�S����6Ti�-�ݷ
M�p�����w븤�ۑ�2}�L���~�v2�8Ȭ�̍��2f�+i'�__R������pVe�$KVKʋ��26�l�� �w�?)�rc�b��k!p�\6�j߸��۴@u�S��G�� �;�d������ޞ�¶�x�M&J% �ŷE�v�ᐫ�F8Np�0��]��I5~��ew// �3���&SJM�+䲿F=%���mg~ѫ���^V��,��iibU&Hh6{y� g��OK��������;��&�:9a�@��d�޴�O�Ef;?*.vsN9{0
Y��m۽&)X�������\`�-�jio���{j6�2�G���������ˋes�έ�$I���C{��p��F�2��j
�,�2�W|�޴�d͉`��X��\��R*�����V�y�g�P2Z�=
�~�A����ο����AW�T$�����á�3�6�;x�k�����z�*�R�Z#Z��6�֐ƞ�^צ�����H��1�hkk��`w����v4Q�����v>��@Lo;��������f^Y^vy�t<q0�qX�<w���F�N,狰%�ΆCQ��5YZ�M�Zr���g�!��}"Uz��w���^�S�I]��C��̖�B&��0:�����wp"�@�aX��i�1��Υ��<�p]٣��N���Fv���M��������GK~�G�b(��f��⢓�bB/ a����@��̎����9)�����I3���M���r:��u91�<�k��_t��Z��VLs�ob�ɸ����<�[��s��J
���k4��"(���費qO<`��w���ÍN�������^����"�������>e��=777�f��������w��	���3���^#���N݄���L�V��W��.}?�{3��`�����UK��0S˛r�`�oT�o����SG=%��d(�3��Wi~�^�g�Y��wZ�U���p}�[��х1�g��0���M�m����U��C�'^QuS�GHW߱��Th~$P�r�?�� u���Emc��W���o�y},���q7�b~QCQ��H�~ʹ���^6�E����{qw+7/�-���'p.!�A����f�X,�u�����.��,k�Q�:]d$R���>���=! �f�L��i�����{���w٦E�8��J+q���Q�qMsg'�8����9Z��||��8�J�i�E��ķ�ݾ��� �q��:ZӺG�=�����T�M�\�.C�C���^wn[��}*�ϊ�Ss��%����fDk�@y�苖f²KE��Tn�˭C),���i��@ū�m��W�U˩?�"���s�Z�Jt6���'r�x_�0���=��s����`�\�D6�vA�XI�n{5x-C~�?ϋ�Rb�ǌ.g,k����4j4���_��ח�;7c����σ�VKe�ζ�����?�tt���)q��\�~p�g��єp懾n�_�mJ�95�ە���S��HM�V��t�G}ek/��9o�VYt���E�g�OL>JZ(k��/��r(��=�Dc´��0��Ĩ��}��{�x^�_]iS� t�2��>���s��δ��@ ��"كB
Y��yW7��S�yA� ��9�'���/_>%W*ⶖ�Ǜ���6�xjf��`��o��l6�^4]9�^+\�y�_�]1z�,���vK-�v{�
�ފ|�.۵}�g?��,v
[7����53T����:����R��V�TSy˹9`��ax�����͵�����=�S|��y)�8�}�c��#�/�y$�3]�o� #��!S��F�ST��l5�n�tn}�#�ӣ�	�V��'���jM�C,|�a1�˗��3�E����jx��`�����%	=!i�<2���3�e!7U_����[�[����|�4A�n�n�г�����L,�"6֙�0�Ρ��-+��Q��1��ə'�W l��F�c������"H+ލ�>��O�&h��������{U�ɕcdh�/�Bx{�/���++���+*�T'���y׉�<�S��o�_���/��{V��F���q����T/�V^�+R�=sTF�Ӥ�F`k��Ĝ�ѿ����kKc�ƿ���{��RL4�'�/��?_y�ús���6)q�L	;��X�1�b���Ntb�1C���j�}8��'J�I2qE�| �sXI�Ÿ�.����t�F&\/�}��¡Y�O�m�fM}�֣�$._�څuR�Sch�]���ȇ&gG�G8P����^������%5:�ݎL�-˿����a��{��l-��.]i
���z�����ӂ�?v��hz	�"��7ݶ�����oj��ظ�s���-��j�Cx��@N|��AP����ނ:�9�i�t��9��ֱ'!?mE{a�"nx�=h22D^�ޑ���y��
�,O-YTʣA�y���*�*�9ttڢ��lJ��*��������x��&�1i�
��FF��ݨQ�0�P���BT�����?k��m|S��Z���n,O�@̎�:e���r'��`�矍 ��"�����Gi����L����}��{��މH�nn���D ���l�,\�-T5�w	-��߮��4
@?�wP�]�^�w�f\���Fn�yd5lb��sѕdOf;����z/2@����"$���+��E�fw"�b�)��Uʃ+E����Z̏Z>A�b���&MH��G������/��d���c��6�Ǫ�+�L�r��}�X�W�mP���$)��g���kL��>��w9z����|2�c����:�[��~N�Q#$�R�s���_ I�F��\}}Z���F�.3,kAO��+q���bئ�W��UR�++��*�Ew|d�x$Y��PҠl�1��3�аT�ض|�̬�x���#������Д�=ZϿ����Rp	-��U-E4S�|J���й�G8����*?\%sr�p�e�R(�������YT��������"`fN��5�( ���9��`���8a��/�W-�P�z����m�ۺ]Hh���0˼���ܓ�Й�����D�ax^g�������q�	\ݛ�O�O�rRb�����
�qlV]SÔĥ��e��"Z�HQ���-�'Ʀ�Avw��/!t����j��/���P̔/R<Z����/999-j�-���ǵQ��h��e�Ζ���Y9��m���{+~���%�一���/�u��*���9�]��I���Kh)��M�=~�i��B�������f0�S�
��ZڵU[N����@�i�p����L��7�;̸E�k�}@ck���K�s so����ʓc�n�.~,��5��{ݣCp�ztEyl�M=s�o��L�-}�/
��jh����l�����Q</��QmO�@��	�(��v�@�t�t��*��<��O�0�]�_�Sε��� �r���]y���fU\��Vbކ�QDHU�nnu�hϺ��ęmk5�seJ�`�¢����)��"�˓]���5���CT�'�����+t�V�]�����.�ʕ)|�2��3A���x��p���Z�v����]�Q�T����{���h��?�����{=S�.�G'�hx��#����Pb_�X&���D�0��	��Q��OD{�8���x����V�!�]��N�\`��g�o�w�'�>W�u�#���<�ݥ=�-�u~G�5&"��Ts6#��UQ�[P��b޸������mj��4$�j��,�������n3��xںm�a���xcٯ�o�����2�g�L�D:�3������?��Yh�5��(�ll��/���.�~��};~�6�(�jX4����� ���%��r��C��J�KP����u�5ʃխ���7���B�v^7&�ƞ�!iׄ;�Xs�� W>P�n���b)R�>sB����mx��b��1=��]p��v�Y>>C���������#����(�y3b���-,!u&�gO����V2��m.����ɪt�e��^���� $�%��+�+�uE:� S�C/
b�ϥC(_���l�� �-�Ż)׾���.���1Ms��)�����J���O��(��Ɠ�3�A����*�.�Z�J�������@4!q�=|}�k;���
>�j�3}�O�Że�=n��⯼��~���� B�N��¤��f�~��ϵ�S��)��<�n���X�B~Wk�J~-{	�޿������w�E���)�==߶&�2_�t>�Jþ-������5�Xw,]���o��P[��6m��������߼E�b|��+��shۍ���MMj"�is� �S����zr�Ն�c@K-�ijXR�g�u�I�qQWc�՛=�YI�A~�>����O8	rHy���X�` �[���g�/��(�6���3\�n�m:k�fj�����Zqv_1o�$O���.�ʓ��7���r+�QM�*R���z�5��"��o�?x'��8P�*��H�j�r�n*$�7Z��z�2�`��%�����bA($�����FZ�u�`��K)��r��8��n�[��I/ml��XX1��{�Z����2�{��_s1��Npw
*��\4W+S�T�������h:����S�ၣ)9���tvt�8#��o��"l�S���T�*4����%����Z�DP"^� �999�!A�e2�+����̓`<e�Nl�h�����h��ih��
�S��Z������x=��(Z
�b*��-�@�[���/��;�3<x������g��ul�V�����t�K�&�Lj��c�r�;�xr�J�Z���n���l���w��e���f�L/U���ym��Z��l�Y"��r��xӅ��:���Z#&�斖ۋ4�	���Jt5�3��fR�E���Re��Bф4�N�_�م�'=1:JC@�C��l�y0D�?��U�X��j����Cq����Y)^�k��Q��=���jqn|�����ұ�rq0�-�Hx�D
Eds=��!d)̦��O6¼��A�y,����w�G���ў�⊥/z<��J�	��aKz)%��b9��u����F�� �T	UJcr)<���pL�}�K1ʱC�u�eSS�c�̗$J��ab��6E=gt�~����P�ji�˖>��
|�H`����3�Y���>ݘ���#��=.`:��~|�MK ����1*B��7�l�ql��	W��A�|fr6��?�g��7?i�&ܜ$����)�9�F��o_���WsnR��sGÆ�����懇unv��U�[��a��h
��4M�L7�Dh���.�����	�|/πsO�V0��y���	��M7��~=}~㧼�C�P -�������ѫ^�H���-`�k��XQ���Ny�W?ܝa��Ǻc���d�lf�"k���;!{9&��b�;��〟�����x3��͞P,E۔���7ڶ�ߌ0S�l������_T����n��(�^���b�o�	�*^O^���J;錶���(w�'��}�
������g.��
�����b�Xv����w��B��[[x�hkkg/���=n�U�un���Дh���@݇�$�:pMK������J�4_̫o��WG(4��nQ��ˈR�tܙTø��2��W;u������l�::?���&\�}ˏ������~�kٌɱA{�[Q�b�$�����%�'��&U����=^ސeB�nU���/1L����r�� �bۻ�x� ��m����S�0Lxہ��c1e�P�y����WZSJb?�����*͈�9�\$eS��s=����m&P��~inn-��l<6�$q�L��B����$9�[����kQM�qv����aBA��l���e��_�Z8���z��ŗ����8��<o� TW[���w���;e���Lcmo_+�rp(���hU4v�d,:"�[?p�&�z�8�H��/�чWr�
���I*�>xz��#+&�o{nI������}:�1]e�W����LN�׸��֩g͜z�ca��ݳf$����3?,�8����Ag7�
�O-�]6�E�HR8~$��M�ȱ�}pG�X/���1g�
����4o��яD��:�}	 jpO{��|�8��1	Z��m~���}�iZkJ���#~���l'~|^>�a���q��	�J�栽 k�ٱΰvlqf#}Bx	/�$=q��fK���/�_�L�)���4�	���Ȥ�5�LNL�]B�{B|�kG[�b��m�l���a�.�9�ڛfBڒ�Y(�������ڐ2ލ!�Z&�gl���+�=h�Ővz�)�M2���d����C<�I�c���0�������pl��OP��,� : �<CBTA�u�;汮q�����{�i�X��bq���Dp���j~~ ��d�c�
��:�Ȣ��Vm��K���0h�_7Z1� d���D�^'�A���ݞ������K��]_͜���
�����t]졓���oF�z��g��DY��C���!�q�$/j�ː��+�������W�UR��R>�ZBB��k��A
$����:�B��+f*a�p��qs5_t�ƛ��׊X@��J�ze�<!O�\��J�%��Wf-I�W��vm	��M��j�j��Ж�k�jVUHP������j���T|gE�u۔F_-��Ls���h,��8����~����Y��A�w�����c\�X]r���[>�iK~�*ꐌ��S��GGF�5�����,}D
�j�xn�-�[Ԙf�4��s�X�&�@/�+��*َ��t�@���Z��rx�W�����w���Dټ!���k$rr�տ?k��[���������a�*o/I�������|E��E�O{k��m&,|�ꆜ��Z�S�կj�"�h_S���Yz־>�x��7Q�g$��G��"�g�bage=t4O��?:b�I��}�������u��t�F>�����|vq�.�vx����&-��3�G(����A�������O���WH�u��#�����T���Mv�N��{�%���|smZ�*ձK�5=Ԏ��R���� �׶)כ�.��ʊ?��3�D�~
�Q9yy�t�<h��c�� ^ʽth1�[[��H1Rqc��+�g�F@�a����/�)�,:�J�zc��o�gaH;�,�|�qצg��E�y<�8�%_�-����c�@�.6������N�i��_�/\�~���)�Q�.��?����'�o&�}q��Z����j1�Q��[�)�e���tE��dk�T��վ��W	u�V�����E&��
��d���x�{��St��ˢ�ߐ�\�J���.��3����Vbo��Qf�)HrN!J�d�U��r��26�w���?�s�!ԒخNܮ��/ƚ*�.0IrW'ŕ��*#�8]T�0_�ܛ���G�9�����]!F�%7��;c/��M�(�'>�c��׫�v.�m�T1\���m����4�ԚO�Өs�+��E7��q15v�<���:�
v��A�n�� ���PLj�\�}�8�գ.�w]ja��I���FWp�m��k���'	wťö����&�ͱEߍ���	�����ߓ�^)���c첨�pi 1��ţ1���)Il�FI:�������7>l�q���g����Y�Z�Pः�y�� F���=8]!|��u�LQwH�~F���omRڰ�A���h{��|�Z/Lg]����?9��p��q�8��n�t)�����4ؕ>��p]SA�^}�$�N�4��X��P���_����֦$�p��,'(�7@Q�����;f�6v��>�E����h.�?{�J�����L\uV�ĺp�^���<�v�����~�j�K�c�PJ�BG�q�'=��ˮ^Q��a���l1��E���������f��^)�A$�=�����bL�g�U�̏�5^<�g�J[�����ru��[�ŧ�����営��ۧ��h�˝��2]pdk��J��;\�����o��r��m����d��H�2�jA4�(%�=��@�,J;���4���n���3��;�l���9��ҙ�G*��y3�}V��ѧ����3�:���Z��U����)��ͪ������_��[�'tb��BN�v^�E?�O��"smfw������Ћ�O8;�������bm)���V��OĿy�ZdN���{f�<�o�l���h�n� �w�@��N�a�����
�S'�+d�_��ń|�?W77PN���� :M�N/��_�%㍑���a/-TI��ЛL�
��(I�3�±�ǌ�8�f�=�˓�랛�w��Qs:��hː����/��Q�0Cz��	�p�`� �/�����V���EP&rꐮ�u�A���w�$��!x��� �1���<t@�{�x�Xh��,���G��o<4ؽL�`�z�6`+�*ANf�1�GJ��t�����b[>k�=ͺ��Y��o~#�D�l��7l�u>UGvNM�&�����l8��EȲ�\�Q�ַc���y\ϩ�>����ֳk=���r�ZU����~�@����0�ٚƦ�-���N1�e��&{��?ZԔޟv0�}X����,��y6����y�Ʒ�����BӜ4��49?�R�����Ƞ�Oi^:��8�^�K>հ���_;�#hŋ��ӅTI�Z��1c��g����c�t��h|ʵ1"��z<xHQ\���B��[��S}cX�ح�lĩ_��7p�6��5%H�w6���VG�kZ:�ew�`���S:&fo@S��%�Y;Ve�t�2���K��:/�Q�!�x��'�h��t��o�0LYbI��z@�\�7\�|��Ro�ؕ���e *���nW��MNN�1�c�-�3�_)i��z�t���W�Q�弱W�'~
��%������	�rɞ���ʭ�Q
��	�sF!�C`����\3#0�J���I�߯�؉3 5�������3.��g����<�B~��:;h�s�S �x��� ��~Y|��7�l��At���o���&���׌$W\�-*���G0H9�L�0}'EY7�����MK�	�_]O��i���>�ʽ*ne"LK�ϴ��w��"9�/V��[nk��!U���R��t�fŋ����$��:�h��;�)��56�C�J�3������y�Vܓ�
�S��%Pf�h��w�V� LÖ��1�hA:�d��z�����T㦚��	��rϘbn�@��׮I��ˇ��b���S��s����I�p�h���\�w˸�_̞�8H��b�/"V��Ւ����2-�MZXz��gΓ���Ʌ����k:�4V �G��[���O2��,�L�E�v��.��3!O @�u69���>�P�,uc���/�6ʶ�mN�1�G"r'sT�=}���7�W���Z�R�0�����d#�Ep�P�R]�q��ؘ|�e���,�Q/��ȹS�:gОP���L��/5��`R�����/�E'm�[T�lN�q���
(�[&�z����<]�@���5k��Z�'�����.j�5�Ώd�.�C�qjS&5B�:�����OM��Е�,�@�}�����R:��e���o���I?���������WIv<ej�]]�:�:５J+�b���,'��QVG���[��aOt�%���~pq�NNm�ו�覤z�T��\�*i�nۘ1����k�L-2�ɵ�)����K�lM��*κ��sq�0�4	����p�K��
��; ��cd]18�Ѻ|��W�
�u�3ǣǂ��r)�W��)A�?UʐC_k^f%�=P"RC���8,�篨��<���H2R���Q��#�LhA�Sr��	�b����͑������:|ӛE�0��2<�����!7���dm.=+�x����4(ߏ��1q���|�����6�]��]A�Co�Ͻ
q�kb>�5��˥�wrk��57��_��ݻ�!ǡ���oMO�Q#�*�QV���ޥG�ǯ��L,��pC���?�&�:�7���]�-Jq����>��tI�_Q��12���D��ӛZc|G�U�r��亞�!���d^�t^%@FП��j
�qǇ!]�燃�3ut
ªb#=�Y^.�����|��gD�S�*1?���C��pwh_��D}��8��a=����S7̈́�;5rH�jNWQ�B"9eKw��f�QK���|m0gЎȬ����v��+e���U_2����~�8:��u��8��K���h�Ȍz�L�Y�Z��7�JNY���vO�=$��NTd`�l�Ł ���3v	���h��dWOݖ&�r�}YG"�Q~����B?�I����V��1�I�.��Ӯ�"�_/^�&���Ť?0��bFQ�W�h߂�a��� P�s���d�9O�y:���U��\��r<1�nB���G���k�N��Һ�O7����[o���[9P�ک7î���O�>C�&�|��PVQ=g-�b�-v�R%���Ҏ'kmh�j���\k�p[zZ�
�������[��)���?(�%ǭ}g��6��ƈ���|�u�h���u&14��ԛ��J1���l�1��������X�YBH�������>J�9�Ȳ��4gŤ��:Q[?�(��A7 5��v��,Nwh��Z���I��u���s˽3D�����A*)�D��*O���d8xQEu�����d��yF�Jy\�c�4M����*L?W��[��	k�~N��G��9�Z-b)mm#u�0[Q�����zܵ(=+W>�t�
�,Lr1#��"�u�������^��FĤ��sudl�6<��лx�_@O!@�R�-�x�*xP8�W�bM��O}�8��؃�ߩvY�_��0#��J�տ���qm{hhE�^� w��r�G�t��a0͔v,�^�H4� ���9[���6��Ǧ�f9	��8*���*��� ��^{�ۄN^��T�'��=��v�]W�p+�Â��֚�s�;��{y{�_���@<��Qv�jf�{�`�ʥ������et9�h�t��$!���+�~�3]�����s��R�b����=p:�J��F��Bv�:<�H�:��7/���Q4l�~�$JM�˘ف�,)��$O^c]>����4�T��
>hi�5|;��X�f"�YN�|~W�֡��uYƨ �����(b Ī{������ r;�{ۀ�m6j��`�YlF%�,�b�p�(A5<��&z5�a��D�����[�*ө�-|�7��m��7�����1dX��r<C��^�^�̝ov1��5vjM�g������2�R&�=����Z�}�K�r^��G<$��3��f��@�>�{�|�k�(V(;�QM�rF���d&���G�TL��R��H��|�F�@ΤŅ�=H,��Xr-x8�����V@~��	n�����!)N'
y'����0X���s�"Ȉ	���y\�\�R%�T��4 ��Ocm�:��V���Cf_dq���qI��<�*���3���,�i�%GMTmzlrYO����4vʯ���uA!9�����E'�����0S���ǔђ��� "��I�k~��yی�q���=�P7�7�r�irt"G]�^�_�\w.��]����[.]o�.XnWBO��Jq0��C5�Gޯ � ����eF�����ڷ�	����X�X�
�?��
!1� �;#�M������z�)�Q_o�:\R�����mǴ��^���)����^#2�G�3e�2-1(���&�X��P������;��Hv��s+R����A$�L���GH{�c���T�H(-��c.�U"JV�g�@j����b���V4�nh7���j���3u�;��Y��H"�m�m���/%�Q5�)%j@�އm1CX�˄�����{Z!�r;�,�<R�J�u8G"���N����B;�J�Lb��1��݈]��zi��(B4w�X;�W�E�L8��+�^Pܕ�y=�Y�����Xu�����&�G������������D�r����=r�Oz�Sr����'d���v�6V�o��λ0�Ү�b���x���ܔ�j���J��]W	�t�i��d���ݵ����[[K�wa΍i�\����&�ԁ�ommŤ�%�������R��W�I��Ϻ`�'�hK8���9�h%{�Z�F��埁p8T�v�����wǯ��NJ������Cz��2�:�fS��t7��Ҏ�&M�M������&��z�n@����F%�^=G����d��/�qz����f"B2��)`עI��p�|+�ҾӸ*`s	�J�Z,ۈ���b���'����I�~o�si�&�y5O��֋�7ú�;��6ˁ��!L��>��y��Ы�a����7\�<*�	���[r�.�=\���Ƞ�M��%Zuu�w�׉��ǐX��T ��+�f_h=��"	���u�i&ⅳ�K�F�m^=�z��s���<Ĵ��~9i�>4����+m��[��AxT�ǂ��aBp��@O//%:��F��?����w���V����$$�r��3x~o`ީ���6���:"������/]Qg���&����Q:�I�����S&2���~�؃����lx�3�I9Pb�m�-P%U�P���)���S+![ZheS>��(�0�y��
� n�t�<)b���l&�P�j�Á[���x��1�:���"�������^�hc�j�>ʄ�#Jh����$���9
�������!���ol��!�v߷Uk6�����:~�&\�H����ۧ k8�V+uWy�S�!�C��o����j4�s��yL���*�2�l<Nj�/y�~�~��9u�|>(��s�i���o��f�
S����^�D�Ӟ�0Lt�����8e�_�N�WR�;$cY�"&�f��G�6��Ӟ��i��j_�CT���EYu����E�#~av��;m"}�T��d}��=,s:=����O�������E)�7�Q��(����V3j���=K�.�b�Al�ثV�5RbV�ګ��~~��y��>�\�^��u��&������ʢ�G�,�W?sK�O���-��.IS�|[b�%�/B-ʦ����j��{����}�|z��~g�ZS���߿�3��"��>�Ipے�h>�*7�(��S�4��*����H�m4��ǆ��%�*��#���e"xͧ=�&A�Ն�t���$߫�m:9�����u���;��<�hZ����S�Snk�w�m�u�#K��R���g=�0�z�s��Ӂ�Mb��|�mEBv���1�,Y�������PKY�ף��Y��-�Ej�Q[��S9u���]�G��Bd:�w�>N#.�k���7A���E�5�?�c}�u�hѳ�y�m=�;80�l���,�/~I��e0���i������������hJ��;F�E3�xD��£�w�W���ණ��7�b��)�ys��?�d[���W���+�s����r�xd�4��ŝhojJ��|0�u�.+���5\��q�!P;�3�j�/^}��5��H���b�6�����˿�]?�}�����Z\/�T7�����ѫGG�"��;��G�뫫�Î������=�g�k���������F�HHɖt9Ox��F,��J��?o�A��^��Thf�4WG��C� �1�=���!p{.��
� )�a��6��̼��d���|����'Qx�-Vw�ؗ�M���4�6��+3ԅ4'#� ��m���G�?p����C{�䍣��6}C_�|��PP`��1��f�j{����$���ai����H��ea��cW�V�G
@^L�bwlҠL<�<�y�B��Ot�Y��i�l÷��f-|�{ը�ѫ�_^A�1	���Ed��5��wh���XZJGT�J�F���i���҂�D�����jt ?�|�֊����u��f23��������y(�$S$;nZ�J� C�ێdǙ�}'��a4�˶"�^���H�S}��5 �"�٨;Q��s��E�3{u�ր���I�r��H.�[�����7$��ɾ ��%�0�w�$Z�S��$W���������Ӱ� �͆s���N�_��wXX��i��bN�잤^�pbt#����{Y=�^��zs�G��x�R%
�AT���Z���[ZC�z�Z����Vƶ��lc�4�2�MZ�mMf�/9�@�����.o�x�ZIPIe�K���i^�$e��n�*��EB�kN<?;�. �L�0.�6��\V�Z�Z���U���/?є>o��aq�}U���󪪌5Ya�Vlz�~���!�o��N�Y������N�J}%-
���S���y|m�y��5��MgX�]"���.��5��٘$(�䕇x��u-ڢ&v&q��4,cn�|f�*��������]9�f��/��?�錄�_�G���wWN۴~�f��� <�o�ϛV7��	W�����XZ�pl�����Η���J]�Ы(�&2s���	pv�%�f��@�Ɨ�]U���&[Kߐ�?�J��m���Ԥ��h�sJ�*�l��6�0]Z5N��"c�6��&����Z�)O��Nss��7�s���>Q/�Y����ꢪ��6�Kz�(�:/0�yu��ګ�ŕ�"��H4��pP����,T��*���P	��������dE|�(_������b�H<��}9IE4P������ĔΌ4���niɍ���.fNs��0��,�R�DQW�<�6+�oI�=�9�2�4<��Oၤ����.�k��%���?�o��ǮX��/Ը����:�E��:$e�^ۖ���*��K���`@,D��'|�h�K����@:A�Ο 'maJ�H�Ⰽ��g\���I�KSHҚԯ�]e��^_���GdCI�e��H��8�\9��ǞH�����* N�D�@F[n4����J �/X��I�4��&l�@h��Òk�H�m֧X�_��kAa�j�������%��ʕ|��h�s��S��ň8������s�#]�O0��>�����CbH��6!��)�G���*��n+�D	w1xNg�w���𕴯��%���v�i[��GN.��@�7��vaA�=T4��bƈ�
�>`e��/h��T����N��d1���<NJ�dڕ��e?�� Hc�'�)/�V��:4�=]��.��/K+ĺ^)�h;.p���'� �,7J�փ�au�/��lj�k� �T�#��j�7W��O�}���K��uR�u��@�w��^M��<ĥsۢ���0�H�VHP'!�-�:���_��/��8��qWy���j����ړ����q%���]�m4eI
ޤ��gU�58�ɐ�M�W,s&��KB���K�(3�<ۙ�)W��l�iX���t�b��3�P����yKg?6J���Iм�L�)��Z!~��Z*S��R�޷7r�X{`��W��z�'�n�������
������ޱ����` ����~���yd�+�BK�ຢ?�_81�����Z-$N�7�sy��$��o�z�?Gw�So)��������@���yB��Kwn�O|O���x3�~�F�m�q}�����bP}�p�NN��o*�1�H߿:�κn����_���׹o��^v{-�aPuo��@�қ�2��MK��V�Z�������D�~V�q����9����Щ�u�Թ����P�>���$*Ȇ_��J�,PBz�9��n\_lp`�.)�ρ ��;U|���S��=��)��v�\������r?l}�^9��*�[�W�AE>�`=#� ��H݌�56�ö�<0�)���\O>���٨�����A ��(�S,J�>���6lp|���=u��q�a�9�b� oa�9zd�q���v��Җ� ��]�p�#��h��u3�q���1����"d��ª#���K+��v1�!y���ӡF����:������"�}��5�fu���MO�Qk����h]�����*֜��|R̃�jt��d7��$��[R�6 �&p$b֟,�o�"}H޼&(���rTB-]�Ғ���T1��Z`��qFr4�?>#�:bpo�������e"�"�N7��F������2�i]PzV�)�����_Z=x�(���%;N�ݘ��,��jl���O�{�q�`c�8ۧ�Q�X4�3�F��0���_�'Kq��"�H�|^�*}��r謺,U�
�́}{M%�G����g����wA�=�������៵	�!���]�g-Ik��v[�����O|MuVMx��v��"Ɯ��B:<������iP���"�sQ�pߖ��]���Să�]��㤉x�d)�V*�
yܳ'u pe����$��j:��M�%6Va��Zl��è������=�����}����B|�(��iX��弦����B(/~Y&U�̡�~��"���y��$:ehZ�'[�P�D�kOYX�=�;�����|���;�z��_hgjײ픒��ΖIvs�k�`���%����s���aT��;��d�f�=A�F������j^�b��`*NttC\������*!*+�7�����-ƫy�a���ǩ�l�j���PԘyS_-CJE�!����?��EO�I��ժ*�pl�6�T	Di� ������T�>U��L�Պ#H��NHֺi�KMϰ�VҸNj:4��B�N�BT�M���wѐ��ꈤ�%�T�H����A�w�e�}�S�2��c���3H��1)�Sg\��B�ڄ��\l̩3��F��Z��9���&ze[I�\����v=cRc'�t�z���>Q�6�@������5�ؒ���N�'߫~�\�!�!���,gD(��|�E2����>\��ki��
��2�-�z�w��5>6&��a�J��c�ʿ�x����~�q?���pLqHȒ�:��a�jm�OӃBZ�d0ϳĐÄ��FG��q�_g�h!������M,!T������Eg��5�f�Щ��>
U+)���O#+%�wIr|�9�čB�܄�;�/
�+���z��)h��z`�p��
W����9}+�~��$;��ţ� S�E���߻*��C,̜�W��^�GkZ��+7k:��� c���jLbY��G��)��p��:Y�5�&�{�y<�R{�k�}�uHl�'�K��MxO�W�����	馯]��7���y�^�wfF�Y"us��0�>MJ
�a�s�KM ��K���C��C�3�J��@efP��*��D���E]����dY��:_g�c�	:��t�<_�=[��:��/�� /��D�'N`����M���^��f��.���8�{��?c4���׭ݥ ζ#^n1�q�+H�km�T��#��W�ٻ����?F�R�/�?��� �����HOZ<���Ӫ9��~�
�/[6��p^��5oN����sIH<V>�R�T��GJ�'Jա�d3��*�6��z�"D~{l\L�d� ��G�1>��2��C�J��H>�������:x���]q�'K���4��\X@,�e���
t����I	Iz�b���O�p
�YV\A�U>7���Yy�F�5��ق�����P�_OH���i(�0�`��M��0.[� �~�ΌM�f�T�˭->��HaJBV]�s�vJ�l������F��<�ǈ�u�1z�1^� � �TT�a.B�{���l�����r;��;�)���02ɼ�b|���`��2��~@`k�=���/Y���Ռ?��j���&� |�ܣ���S6��j�1c(uA���C��<�ȸ[}��j��Lu��	�_���6K��:OII	:8���kk��8�̾[p�jX��#
���2�$�SAyy�}�]u��|,��	%�s�e���\W���V�>��M��4�mڃL��yuˍc����N��y�g��I�>�7u/�	h B秦�-
36ӏ���v˰p&��#����������xx�t���s���'��w���3���y�cӬs�j�$�[QsH2\�������2����A�dHl���k��h��!P��So����>�{__Z�w�l�n)�!�8�>^�αy��ÑA'�-J���Yf)X<r��9v,}A���Nӂ�U��K_�Cl����*��fŻ�e�K�j���xG:�a��`W�,	Y�+q���Q3]�D��)ʜ��uy�A��y
�{��x�M�0=���L�l��dST#ܾ:�r*c�>`��5ɢ�ݩ�@%�c�v��i����nrc���ʓD
Ww[���-�L�!�r��V:|��p������5F��k�D��,�B�v�]���wy}q��2�-��J999M����j�.˝��u�ר���XX�_�|ˌi_�'���%�� K���>klT�a���t�����������W�|�rQ��0![���|..	�$%	8�S�{߻������2��eB6�%b9R�xřɘ�9�Ad.��o����%���$~QcS.�B�Y.S��vR�<�:0ːؖk��1���d�� �#Y�\�Vc�,4v���j|��k���dם�?������yܶG?�f=#pku����4���W���ހ�WAF�������a��j� lۋ�S
1���r
�`������D5��d}�)gA�y_J-+w>| `@�j��f�0I��]A���\���ő
3'c��뀝oX;;�U�Ƽ~$Z��V��������Ŏ��ƣaǟx��;"����>VU���6����.�a@�w�u�.)nc6�?��z�w}����.AݛY�������o���s��R�<�h¾��˶�ΫM����~x��[���������Ϳ7��;Η6Ro���.8��߼n�|��0hW/��Y�%Y�Od���pul�>I���cY��p��_�>�ٕ����ci���w]�t��M�TV��]���{Z�b��.N0�@���T��;�����f�NM����e��iO�j!(��3�_G-����JK�V�E0�<*J��[W�5xS5�Է�M|��_P��^��Ƭ�.�[���c��SA4J�@NIŕ3��Y
�Ct��IV�W�B�T?-�r��f?��2�(İ?P�Q���HV�O<��iDfE��I|G!7⣛M�:�*&'�%�<Z����o> ]C���U=�ʗL�{�F��Y�:`?i5�n�Գ�=,]�҄%�������c��ߒ߯~��lGVⱗ �w���K�Y������Y�m��A��>0���W�-O�B9�����%u�ȾP2TM@��q$��s��4�i�t�~/#�0���=θ:>@r����$�قV�.$l�����+Rī7������|?�$�ѕ�7媽������l��hn�{�-n3�#�I�C����ښC��3!�"��1�b7����i�W�D���~q`6�I�e��q2�nw�n�-z&��Rx�7���ROO�"p��72��9����R&�9�����۶-��5��&y�`0����1��aR�{�	�����/!�Z�<re@%���
Q��5N$?9����=�Ɇ�Y�9�U�RSXH(��,��7S�H��R�t��*�m�SS^~u�O����c)v��3��"���y��8h��ܜo���4����K:���B��s�Y�32���aG����y��<��{<�<��������{aGõ�pF��@9��j���n�tra(���.����b�ǲ�V�߿EuF������������
��B��!g�����W_J���� ֈKV���:0"<5�(��\RN�+���Y*���D~�����ۇ�j|,o�:���1Bl���N�W3+R�����=��_E�	�0�'�  �c����R���wƖQ
Y�D.h+%�Z+r��e��xfm�3�M�]XC����՚�d�[���d�~�A8a�.s8ngУp߁�@3�������ҿ��{ g UH���|y�6����L��Q��x`���d�r�S�$��>� hv�V�[,�y�����;־Z:��o�0|�9K�+���f(¬W��M|�W�UꢷL��y鮴ؔ�V�>P��FT8[e��g�b����
r�"�wY�='��ʜ��rE��-���Q2i`+�B��H��ۢL�-64���I�a1aPaE��h�����E��}�����ğ���c�p>o�տ-~�l|�SM��k�d�)n$���h�m�B�/�k9Э��yT[w[���� ��5����+i24m��'Eo9*S����`t���Z�9z<�bU���^��	����Z~_w+1����9�r�p��}������T��Z�Ƿ��LSp�:#���� ��c���&�D+���U�u�m�����q�1��O�O5��ִ�N�S�Q���4uh�<˙k���̾�T�ۿ-��ʝ��ks�o�7U�	U.�K-����"��A:�|S�P���7K�OZ��5j��(�g�ى*6�6/V�86���[�ˍ����nI)�@�9�қ�E��+�45\5��ν�~"P��c�0x׶�r'I�߆,G�/�ߏu�|"G��nq�R�[,�<�k[��)��@����p" �L��2���b�����41�ӗ���K�9� �\�m�߀���>.���0CA��>p�����K�+�V썡!m��A^�WT�T�w������o=~��A�73�e�SGR��%ۛl')-~m��,~��y���Q�+�(���t�4���w����z���P��6_��Ii�.;	��=���C�
W�L�F�^�(�|)heF���Xe�ł �6��d�U�	��I�r{g�oUc�_]�hHGϹ���^��hČ?ئ���ϫ��d�~���>Ӣ���'�7���%� ��MکŸK^⾉OA>���M?���D��I�y��	�o>y~��O_?���!�ЮԐ$j+Ob�~������b˸���\~��<vS�e�:�ب@��;�]{k��#�����S�X;����ؗ�8+�7�Z��췐�^����7D�xV����r$�=|��|8��Qm(�>n��o�ؙHUb���j�]�%�»�_rΔ���;ci
��~����Sx*��+u'�c�"� ��,�LV} �ʀ6�Q+W �1-f�飤�[��i?k��8�(�Yq[;�uп�J�v
1�(z�+���Sv���vR�n�)��F�Q�	̢!�85i��W|Iа�澊��,��o�y�����,dv�QW�|��bĲX��E�R.=�9�ț+���>�}{9�'�56%�P�b�<�s�;0R�ǘ�������κU�j����*dmV�g���ѷ�C���_�;-��>%��.��ѵiL�7�*d����rn�%�}ό��
��Q�$������-�g+ywz�L|n�cQ[- �u��Wa�_���c]�y�ˆ�QnLq}�+��w���X��o�ԧ��<^y��d����^p�� �;��l�3�>���o?6[��Κez6�|^1�U.��/���B'9K��7�ۘ�M�o�AQ�G��%�E���o�6�r����妶׿{w�0^�w��I{���<���	�.���j���]-vn��#v�<F�VtNv��t�܋�yӒ�"gt�K��q)��xB�x /Ťd�"�{��!EH����)�@M�9[�o�w�������&0�"�<�ݿ�GT��2\Z3����������3&#IR�U��%w�9����x���������Đ���望d�$+�K���)�;:/P�9)j��Jq="�U���K�YQ:��/��������"cÝ+fl�C�g���p��U��{y_<۶��%�L���u��R��5V}�o��x��qw��-B�%u��"�M`��,�|H��9���(��zIq���O� ʔ�I=���2u������ �Ùf*-;�p�ћ��Z1I�P�,�`j��3e�!xv��vܿ�E)F��dA��g
��B/W�:�w�CԵ	�/�P8�*�g��@�<�b.ٱ�m��Bm��w�Um��P����rz�$�r��#��(k}��c�@ �Aڕ:�|�\��e��Εm,��zz�{G�7����7�����Ac�R&��Łe�Kj���(��)�����x�����~�'�|!d�Ac���ŀ���i/���D�d<۲{jɮ�ż���OB����U�	���'�"���'N>yZ�X�k��x��`f�1�Ev��]�n��g?2ML�4���`}i��u(�A����Y��@����Vf�E��,���*o�q��'KA)�,�&�����֍�������?iw34,X i�#9��I7�f��t��<�.���n��͓�K�����i�q�������[H������.�}����+w�j1t�]�f�q���i\~?�o`蠟(��|��h	��S�^�CW�'"4��D l���]P�������hS^���p��Ɍh�~�}���He��z�MWEz�&W�A"0k����㉙p8�F �
|�Tr�4Q9aO��۠ 9����F�YQqϷ�ojo�3�\_\�7$��嘳,�<8�fn����*O������ݻ�+��L�'��w��1Xo�{�L���Sd0��]��6;�{^�ţ�]���+�����h��9"K!�(�!.��q#�Ɛ���Dʢ�(�1dƾ�`"�R�=�l�Un2oPt%zI���.����h.��[�I��Կ��H(�zV<��Ä���vX2��jEE�7��y�ܨ.��߮�Ҙ��ϛw�z"4��������B�l�_��}�I)�(}���G�JIN��Z��6��~RV
#a��~��8���瑴ZC��-���ݫ"����+�C�����LE[<Et{����c�����w�̍�C��w����ܒf���i9�U�0�q�k�w�s?��--R��C��������k�&T8�գ���0`#�K��S����D	�� �Α�[f8ݖof[7�㭷��������Z<2�H 	~)�=0K��? ]�-��F��yCi))o�|e�o�.w����ߎC�%Z�����L��pie|�B�
���e�� m3:0�l���t�n�Y�s�`B Y�V�e�s~�����oC��3��i}�����~�QӮ�'��xZ�l���9i�;`N����ü�V%.~lXܫ�b�W6����ߎm�?{�m|�8������M�$��O�|�WB����!�Y[��z��D9[�
hf�<��4F�E��"���lP��'�NǞ�x�G�V=42��N�he}%�;�v�~�*zC�uy�P/E &���j<h�q��Gyh�M�dÂj��|2
�D�U&4�
�U%�!w�Up�7���mj�-�k��#�@#�*ugn���ö4z!�5����̵� g&M��py풯��0ΝH}��͉���D,�O���X�˖�M;Ow�8���]D��- �6/:�6a�%ƍ���y�\��ۖ>x�e�����JS��O��q" [F��FI��U�c�z؜D�]|Y�|��Yn�W�,M��£�'��!����ZQ�uj�Q�D�����h&`�SZ�d���i��#�8,�H��+��]=���L��}"��,�qr�e ����[xu�,~���(���Կ�m3�P#m$嫿�<x�Q,�Q�6�4I����Ԝ�|���$v��b9�#�Y�g��kĦ�:�-G�Ш�x.�a��8|Ԏ�%}��Y�E,[�5�%y���ʇ/s)��y��4-y�"��<|u�ׄƹa;B������&����s�O��s�� W�Z&���$�	�o��]բ�+�U���e����c�<G��aE����p-�x$>u��i`FGyA�+%��xϩ�~��wa���rh�1\�*��\���CLDoj�36�
\z���p^_ tm��c�"���FtYHwҏŤ� ���q�&SĲ!�Tl� f�`4�4����KW�"���,���/`Ttn?0SM#��J�B��B�2��
7E
������Tq���L��a�>fA��/���B���
E�J�Q�G�S5q`w����Aj����NOf�>ʐ��������XUoI�p�e!"T�2���j��{�0h���ۀ�c㥂>���7&���s}���s)4��%D��X�ީ�U0�E���5ş��)L����߱��o�����)�!������a�<E�ϒ�w��Ή�{��gG)y{Mqc��M��_h	w�����O@L����AీV�Fz���V���T<O�V���/��hP�����L�#��A��6�%;n������Ck*�-�� 彗�L��OYS+�b9�D�Sp�΁�U���S��zK�,S�4{�s}L�����ˢՋ��{WS��Qmm2���,��6Yii�x-2=N�,,���I%O.����1�t5�&�B�i�2���f%ȴ�)����=�*�1-�AElX�[Dz8���-W�՘�>4�њL�},Od����X��'
��SP�a�yX��i����l���f����dS?���7^�L��}!p�o�{��T����m�+�(�~Px���))~K>�+iI��trҐB�A��à�/;^�-�ȯ&��$�V�1��s ����f�N��Z�K��A�m�X���E-l�Ʃ���f;<���`�T�U���=>��$ޙQ�g�NJ��R�I���"��?j���?�]���`,%K���y���ED����2TgYC}�x�/�><H�������4���L|����0ep��W�7��a���+d��Nw�T�`��;	�Ⱦ���9���x�@x��0˭�{�, �Q�y�����E{�Fi��[�u��~�X��MZ���zG����s�V/;V..r�|��G����>#�?e�ҳkP��urc�x{>�|���0f7��ojJ��%b+�h���D#�^�i�*{�&�C=�6(n�R��U%%R^�C�\y������n�ړ!����w���8��	�`�,���$<1O��*�A^:�0��ڗYyG�os��<�5�Z#�v����6Wtƕ�<�Q�����)$�o�����=z��U��j��/3i�	��W�_���0��/�K󴠹�j0�"ސ�68�ϫ �̲U��P���v����v�/���Ǯ��+��S�V���E�Wr;�y��]'����͍M"��x	�c���9��z���ʛ$!�z��`Ʒ�]����8%|ᆓ�ˀ��z����!�ǂ�>!��Wa���S\�:�������+��t����-���P�V<�\�bU���a�k�u��1#+�1��'�(��+���,A�`z<\3hl�����Fp�-��]r�������Q��2{����#/J��B}��!D����lN�]�;C29�%��TL�BŜe��4
���������}�X09�N������ܟ?ȯ.m�85Uϸ����a����Kr����y���=��u��Q�Z�	�"�7���w��ሐ�&A.�*dbr��;���r����(��>{7�[��8��I[â{N2OL���:�L�O�԰`�Zh��8O���6kL�~y;�X]'��T��-���DH�C.C����C��-K���U׃��=J,_�.����7M�]V:�'����7!"9m©�~�L-Z�o��?�y�3!�q|����O��9m�pX�A7C��$o M���_�և��P�\���*8���>���R�B�	��� G�1�T���v����~�B�s���K)0օ#{��H^��'�AU�*aF�t��'<��O�?ckEM_�۫D�m�6�xU��ufN��
"�َ��Oz���@��gٲrBO�:��d���>(Ո.�!p��&0�4�H�;�1��<��p^f0nR)��M�I\.�xǻ]�	CNB[�=���E����|P�����>ʋ-���4�r�~�t�|Fifr�3/���*~��_��k��y�1�ٺ��j�۬�k���}j+ª3(�<ԦޛHH�#��{���rՁr-@s��l���i�ʵ<����w���[�L�q}���HJ�ä��P�MVw���O����[0F�Y��a6�f)4�/m�I���\��TDg�8�|�؟�]i�x���1�e���j��cğ�7�ϯbE"���=}B�ᨲ5pcf�]�y�����A�!�w���O�2!�L������ɉ*�Z�OZ�S_?U���@��9�y���6-�������iޞ@�vF���pQF�L��@"�;F]n���<�'{Yg�/��<J��z�Y��X�Xо%��"��W�/��ף���QgU�R�@O���D$W�/=���+��V�=e������# e%A�q�SG�����H��rt�_���h�rE�k�KU��u�r�{!}�[|َ��)߱H#n�9�yXI"��k�lM]${I��?��OK�K��3�ݹ�j�Y9N�tޮ��Ր�~�������Z��Wn�VI���	��k4yBU�C;ɟڲ&I�4��a��ik
t����<��v��z-~�k�1����с��~�������wd�K��t��!3�$v�
���SW����T*��y�\�#� �Y�t�T�N�W�hm=���3�"�{��_�}&�sP�N�N�imcspq�Z��F�7m��}�3uʒq��S�U�*|�*|�%��l+p���b����Q�U�_氪�;����ZONT}"�z��90�e�����X�o�*���<� �w	G��}���5�2����q6k
�6�5c����ѻo6�5�_Z����r��O���v͖O�5��j|`k+c"���;�7�A�&_K���-�r��}���1A6������1J� ��\o�F�S�p�	 ��Q���4�؞�y�KS�M�2XB�x��b(��g�&!�{����ոz�s��ѱh���i�v�r�"<+�Ѳf���x>Z��������eH�h^G�߀�ok�װE����p���MN>>�Jeo�������w��n�N�m;wڻ�o�~���V��g�Y(`�+����DMC�/|�Lq�\��v��蔽My�5s2{��0� ���v��.�C�͑�_M믷�A�w�� �ٙMY����^]�wD8G�;�r&��uZ:_��ے������7����M�Ȁ�Eh��݇\t�� 
!
 mR㌞�ս~�a�[NX��KH�q����rň_K�R(�����V���"#Az��|PJ47y5>c�zc���/�߲k�^ދ�C�tɗ����_��4qʥБBx�������CpƦ\kZ��㮍����7Mub�E����>���h�9���8��c�П8e�����|�YE��{��*��^~���9�r'/)�!l��q0��fhF��k�y3��H{���:2���OzШ\0b�Et2g|s�$	8τ��w��O�E�y�`$J���` �Dv�����#+d�A�_H�W��k�Q�I�9�������lt�m�����Rkj��mV���� 's|����_τ�c#�8�XW���jn^(u__w\H���߽A���C�⾤����Ĵy?��@t�Ϊ6��_��;Γ���'¢_֨&���efJ���~�i�n�<<L�#���%(+�2I��*�^��h���]��5��Ϡ^�tl�A��n��pB��͌�5OPg-P4�>P7�N��Ko��c9w�?v�4�iz����Q���p�7��>�ⳄU륛�>r�\7ڐ	J^�5s�>X���;��;���g�m��z������*a؝0黖�%.�)�D��N��-�q���zu��-�1r��`F�v8�-+��U����0��{�������?�Ǘ���G����dueN�����l�`Z.�G�a�e��oI��j�s��W5�����x�qR��eR�EW�0}PʃjJd��x���Ď��-,��[1��)DTu���dR�{�qkk`��ۻ�� �jmv���g͜f�3�fOc�_� D�>��UڤOn��������c�f��?�j��9c�h�ho��R{pɣ
4�9v^���5kyݱǳu��m�"BVΜ�*  �b�4�7�VB�Py:P�8���3��0��3d���{~��p����C�	k���������^�Z;�ɮ��,�O��
=<΅�o�N7f� ��>�I�f�6�d?��D���q 2-@�|�)ur�I����ՕƗ���a�<5 f�Z�F�����{()SV'�ch�ⓒڈ��$^��ڦ�5�}*m��k�ݮ����͖�;�ֲ��;w��L�^c�!��g����B�!\x���H�����%5I]\{1�4�rQE ��_&��тe��2��(|5��kbdɔmC)�<���!`s��To���;8�U*�x)+'OM ����s����njQ��|��d�u�7�����~�[&�9t��Yh��r�#�~���l��w4c���;fo�Z��>��Z|���-|h�����y��N��nǾ6&9)镵ٲ�Sy�4x�]z��(}����]��ܥ2�?�uZ�<�Zۊ)�I/�.�K"���, ��0�[p�X۩��b��r����}Mv�!p+��=?��� �����EرX��P/~-'�Y��v�u.���5�@
5�����q��j�hu��PH���F^��P���{w�v>��R*h`��)�^�e�I���΂>,vؑ#�U%�?$��ꝋ��Ene�o$*S����|�cfR�~,�lJ���S�++�PR�m�UH���}�%a[���?p�I���ͻ��%���a! �k =$�]�$�R�!qem���7���B�j��w��V�%'
��\�h
		��+b\8�� ;|{�pW�K��rP�S���g�F�E���ݤ��x��&A�~�����ͺ���ȃ���D��9�¯��4�s����+���˝t4/:��X�Ӫ���G�D��lS>I��!tS��{F��e7�o��)~�������à�c̱전�.~�&�g�&�s�$B���;�;i	�2����Kc���~�UΗ�f7u�]�F�N�(��X�s�4-�s�J�������1l?T�����bB��4�Y��#�0���3�e	�'����d�J���[J������T�;�4��qR7.��T1ضa+y;�� ����]�ͦHCq��<�^�����Д���xjReFe��Z=�=��0zA���E�����W.yyÎ�����ރ�3t��6�Me$���*��
]�:�E3b��.l�}LX�Q	(%�j�N��O"�R�)�	��e�5׶�p�k
>+쳹�*����k��H:��o��q���ۛ��0�4u����6�Sd�wi�,@R&�����z��I���nЧ�.cV�|�����4и���I��qt�qM�]G	)i		%� AB:'9:��KiF)�Ȁ!���? 0�v��g>��bo����9������9E�Bmޑ�-Gt[�H����9���O�N:Ml@�-\Q�}uny%��T-�|������>��e/^8y�>�٠�޽���c~�Fmk�h��$�_�a /��Z�����;�I��'$f������8���DK�X�Z��f�y��ӷ�K�e[\0���	�GՙƯ�1���������r���z�����;h�.8_��"�G;�QNy���=}�>
aHU�����S������FC"����W�t�F��Hw��K��7�V�G���Lޒ�Nϒ��uo�*g�E?t�W�Z
|�6��}�N5���{�Xd�� ���-qc��bd.�KZ���~�N��7	�-�k2�ށgjzb�J..�H��i�F@Yٟ~5��A�++��A��^*󆡇f�osv�x<���Sܝ�Zwb�xfwv 	#O�������+6Ȱ��(,P��t��!	1�������3>j�����$YNa��75�����{���:y[�d�Oƃ��V�ϕA�����HU�H��zп�f� ���]����@6o�t�����:�"�k	�z�w���9h���1�������k����� e�J]�%Ղ��e"��5�����/ a�.����R�	�'������[r���6�P�����Ӄ�T��*�3��|�!����9zD6�a!{���S��6�;���܌��?��a�O�~A¶$�����@h]�[�h���x�z����f*�JI��n���VY�����
~� !�a���< _�W�9������3��$sjL�wL�H�$,5mpE6~�{�V�~��nB=क़6 @�ï��B����3�#<��Co�#`B�-p���ʠ0Wń9]�|������A0��.�ը��V�A�c���a�7�0�Ӫh�s�/,���F�^8�r�Q�jA�t�\n�B�����m��� Y
���
S�j)���QF��2����;�gr�+
W����U��}�Y,C��ԟ��,H�i���y��/�nEE,&���	(�ل1��F�R�zUv7��Ҏ�
Ҹk�� ޭ�:�x?��V)�K*�'O�gʝ`��jW�Y�3M����gp�eɢ�2~�ۯAj�6sv|jV�]� � ������Ӧ 02�O��C��}�K���ƽ՞$v#�ԏ^��N�X�P���$��&�
R���܁�ߧ�-�v�M�okF";������[#A8��:0SH�d�+W��~�Ȍ��׳bA���?O���66H����H�n��]-���(�5�/�Q8�$UM���,{�� ��0i�05N:}��o>�O�P�瘚��?V�%<�X�C'5^�Q�i�{֧0��Q�lϕ�,�t��@ ;���j.��/<>,�,��@kZ5�������K��>�ǉUl:e<�ݨ����G�F���,:����O>��1�Al:��*& �N>xe$=�,^��E�� �`���������f9Z��~Q5w��_Cy�<��R0��p
.pU�e8@�W�F[����Dx�"�1Û��h�il-���^݀�Η^Y�6Jp�g�1���qrxm}[��������<����]m��H����X�w����2}^D�g�2��`�G���ȟ������������.#���\1�{a��MAyֹ���������V-�#�{vv\wYw�~�{�?&�,��t�ikkK��f�&�^�Ϧsн'��� ��8�
%.�0ܬ���#v��{jui���m�W��M��G~�����沞���[5�h�i�������-��S�pvidG�2��}]�Ӭ`Y,�yS]�:�hWS?�:S�����)����w���m�h#^KLJW��%�E����gݔT?�r~����k�B7����+�/</NdJn	���	6m��
��P��)���h�h�H_*���?�۾1�q��:u��ؖ:�۴I'���-AԽr3o�N��a�ͧD�C;�� cc���M����CK����}�22�	{�������է��֐Pt���_xU3���caf-zn�%],����r�"VI�Mn�?߂�Y#�ZD��������^�/to��!��*�i���o<E~�§1u<n�;]g��b��4����:L���r��%p��R��+�񤳹2�(�=�j�^��I����	�Уz������uU9}J_;<��c�ݏ��ݢn��0����N+�>���
�.�ðT���x	�:K��QS���k����f�H��m�]q���+k�`���9!Rh(��UBb�I�$#I�4�l��^8?����0.��%H�hYH��7��N�]iߔ3���.�c�6�?IB�/SJ3n849�bH�j]����]�1m.k^Mމ[��r��v6�x:�86f+��F��&��i�����k��Az�-�����E�L��IE�()�Ӏ�u���@���&��r��t�]\d�Ń� �m;U�i���S0�%yH��Ywubּ{5C�q��������tq����|�Yj}K�('�J5�nuf�����:���S����o|�̘���jtb��K��e��':sK0�T��l)��ɚƫIG�8������ev�z��N�u��0�D��`�*������V��zF���ز	�a�>g�z���	�T��9��&R�	�W�;;�SJ�ϫn���,z��]vu9e��}W�g�x���:[�q#�X����Z���q2?�F��8���|aAH�G5�}8C��*�����)�I6+�0�.�W�5���#�@K.�rG-%���5���s.k�.re濿>L�O���>�����������z��>b�x\t�f���e��I����Pďl1:�{�6��f�X�S\����չ���C��i�O��Ƌ��%c'e1�)�zoI��IP��&���bK��4A��C{�d��C|�v�RN�'lؗ��-�I�(�8���}��������)U�e���?,]��-FG��bl�и�;�����h��$��Y��U�4�E���>'�K㼻�V��y�|�)�{a��:K[S�w�=���zn�{�ϛ	Ke�pq��9+���HB'�|���.��`�f��A}�7����/hv�b��zڏ����}�u[&�z�.��D��B5�,:��t�Y�tF�g)�.+u�ٔb9�Z�X �r��̀�����I6��Ee��Ok� ���,�&b���uګw�T����VVҩ>_�Zfp�oD���J��O�*�^�3o����k��!�G,�),�������E;�-��@9�4��1:��{0���y��f^������� �%�|k��i���c�.�<ݝ~#o'��d`��W�zrqv��{2Ig1��1s�ȬJ��忼s.M�6����f"_�&����3)*�b�4?��a�{O�,�p�7*jѩ}�,U��4ձ;7�x-,O�����c��}��c#g6Ծ{�L����4�����i���[�, ����s��p�]����^&�؛���eՈ�{~ގCb�����h4:�i[����)081/*FA�'Ӊ��KWՇYnU�$1P�Ɇ-L�2SPP�H�_�Jr����@p���V�@�F�&OC�l3[DY6�'��܇<4����^?�IX�Uy��}�Y���*y���K��-�0K2!�,gG�[��K?r�1i?0�)�5�O�'�@k9;F�E�|�-��.�Y��\�f�wA^H��?���]�h�jW�s�s�T�O�G���;�hC��uc<�q%��G����R���qP��OO� �?T T!@D83\��l��T��d]��ɟ�5��t�&�j�Q�o*N��P�|�J�e�����]���qʏm��Ղ��|��W�]�th2�i�|F����w�\r�껗�^����Q&���Nw�ܜ>jJԣ���P�*�S�S���/��Ah5ˮ���1;1-V�i�K.�>g�X���\��eNe�����$�<t,<౴��b�\@@�/�/�1�;����jY4���=ߋJ=;@֭K7H�n�\ܜ���bZ}k��_SǾ���5ET���M�z\d���-|�=���Ԍ���P����g��������7��ϡ���+D�ʽj��!}$��#�ɏ���
�O����i�������&��w�"ʼ�5���9��>*�插���������-ONhǟl��S�SZ�,+5�$S�r����yf��>?��aQ�c#��⃴��.�E�"`)�:g{���*�i2�偤�κ�F+����n��5^��su�ݳ|ssU�W������G��.�ن�m��Dq�JGF����_,�q��kw���U�o��߂.c񌗅��#l��x��[ƾ���15W��Hc�d
}���s=HE.a�U|�B��=B ˓AR7��"m�Δ�ݡ�U�װPyN��7�l�a��k+�OY��
��K�\��
�0ggӍ�yle*�Gg�zw�}��%j�׫*_���?^>��2��^X�G��<(kq/y���M���;q��^�}s�����ۖ�\amR�nB-�Ka�oeHߨU��~B('!�J�666��&��e�"�j�9���vh�U"X����\1���N���;�}��@� �T� ��ܷ?���/���e�lp}�}л��I1��b��`E�Z�{���L����pMa��7W�z��g{��kk3�Z\0c�� �u���S���m�_8|�l|"Ef�d3$�+��ψR3��8B�O>��e`�Jmrle�̳�9���D%�$S���nA	[%Y&t����a"% clN�lY��c\�),2�'I�nk�)�^}Ǟ��=���gm�(Z���e�Ru�*1rʣ.�EzX:sum�P	�y`zחNv�����z
�x��^����HKeV��v�cK�&D2e?4u�6�ϡ>��'�>aԦ��c"��X	�x�v/j><Ή�y�#�N���� ����&�Ž�[��N*:���I(ޠ���� �V��fIΑ͹���3(H�����+�g7l���:�}�EUu6
9<|�c�2�T��P��$�?�'\ ��z1}g��wr�cG����>�Y��wT�?��M�
_�g����A��_�n��]�O�->}�>�#�c��&hԎ==�dR�v��,i��gq�/L�XG�6E��t��lu���N�����+��V[G�����A�Xkϰ�Aw��}�\�\j9����rP(�9mzrk��YW)Y٥�M2d�٠`D�� ���űˠ.��g{�m��	ĝ�L� D/�-e�  ���X����{�s��_�:ي��F��<'��v���Gy�f��qI�����@72�*}��0vA���7fԧ����D�<�"!�6�����'�$��H���^���d��gQZ�oω�;��KHi#�T#V��@�D
�#���sQ���O�����O�����g#@��۵��`����I�ŀ6�ɤh��>���W�2uA���ϋ�Etb����,?��ى���������?�,�ZJ�������g+��8��a�|�ADx�0��n3vؗ]���,�Y�������=_N?$��� �P�h۷6�mk�Ҍ���\�6ֈ�gq��5�Q�R���C���p�*��]�i~sQi�'�]X�3��
���i"��+� ��%���S��.��YY*���҇�~*�e��Ayݸ˂�9�wb��7��^���)���V<�����ǾԐ��C`����9���]Մ�/�0���� �GjB�ǐ��OS���߶2�r�g�EEE�<�����"|=O���e܄/]\���YA��:���\����ң1���T"	0;Y;���\�� ���)�������U�����8���Da*%�/�������i�֤�8g���,���D��9��2)Ul�d�W��p^@������ &{!y���H������*J�u�s�E[3�Y�d�x)���fO���6��Ӣ���g��'�rrB������aׇGXְ+J��_k��A��5��x�'���Mw�N�ErX� W�kV֘�� C�����`�rNz:Q��t6�	�W���
y��,0y�X>�^$�����n�	�KKQ^��v8��S�e��S\�)> ��$�+de?'�q �L���~ޏ��n*����2}ɐ|�^��L��Ƀo	uh߫�6�͚�Q@��=?�c Ih�(2'�Gp]��"l�N-U���!�2?ӭ�_C!�¼�]��k��t�hcht�Q��]�_���d��`^f�}���K���2�&�繬�NAA/�=��b5I���zs@� TѤ��ԍ�OhR���a�
���n�\2=%�]k�@H���g��Ko���?���	��)���pj%�3���4*����V�@�<�|A�<�nf��ˠ���ppf�˃��;?��fw��`�2���?�,�fzx�\'�����Y��KA��cNQ_�����áe  0��ՅZ<u��d:�����5�Ix�v��1�
W��بb�hi`Ԅ�$�HC"n�L�5-��
��k���m���✨9�<�?���C��;���=&��TIa���[�r��EW(^�W���AJW/�{��f]��-is/-�"n�o�Q��kރ�D�����Q��_�7�u��k�dQasU���,�v�+3@��E���×y�t�al/�\�,Ç��<�t1}�969��^_)�u�^�R㹦���	�b5��[������F��Z5I)�jto�\ա?�p�CF�I�k=\�s�xc��鲘4�3��g\M���:�o�T�oH o�}]��$�N�(%h٭?b3!��j�k�ѿnx���(���PON)(�Ikп<�Q���Y��M9[��W�O�|/Q� ���P�@���?jm����w�Y8�ޢo�M�
��&[�ɮ�K,nH񕤑��[����'�˨n���ߩ��a[W��HRӡ��)	#�q8�w�H(��c��a��$�K�d���2���m�H��*�n���K[Ψ�]1'uph$�}ga<���2���e�\�K?sݓe�$���/�߅�s�W-�0��ƌ� �o���Hm��Z�̸��n��H�_L]�J� K��.�Q�B�MI(��b�K�ڥ�����Z喟X@=69�w2C���!l�#�y^�$k�9_�?�dZ��mM��,��D{������i��[f��DH3J��Lq2�jy�L���C����������j7~�-����`�
��t�� �;�K��.��v�3��'���([3��y�[iWμ���J�p8����n~���R	aߔs��Ѵ�O͒�꧸���P1�/��'����T��ʐ��Ts�Pt����N^8xyݒ��ZZ����^x:'-��΍\w8�|..�`-�2�Y|����ʇ�s�;�e$O��oj����~+q�t��v�^�>9Jyx�98���.t����.�K�z9�tC&�项P\���짷�0��WfD4����U,XH�J��:?�B��c�p�y� M�w���@Blk�A���8̶�!�!G�E��mT�p��[����Q@�W����)�i�	:0'}��7�O �fnN�(m���d�ԗ>�ZxG��Ӭxi��t��.��M[}�����<��-C���܏hc�w�5�gCkU.ۓ���?������]���A�����D��!fYU����q��S-ҟ��Q�$n/n]�T�~�;ٮy �� W؉wo���P����B{�
���a���[�1q>-��FU��ͪc-o�u���5F\�w]YL�q�x[ՠ]L��dG~��ۋ_=�cBM���S���_h���/�d���H�^�JQ)6�Y�R��Jp�c�pL(��x��?H��2z;S��3 �}n�P�v��}Y��@g�t<��|ݧ�Zz�(ʑ�8��+���^/��=8�d��9.����p��*$S�r04�h�"J�2�j3��+�7�ɜv�Y�a��Y�&�֡N6��Fe�h��&�����p
N�����9 �9�޶���TO�.E-���؋��;:���"�)��4l��z��}����1nǢ[�L#������&e6B=�׸���A�' ���Ч��|I��_k�~�X_��U�9��8�F鐖ŷz,L�iEպ;�~W����r=��2@?�@�U��󿨂��IР�}sJ�$C����W��<(�~%����
��Lv�(��/��b��]/�#.�o�p�Q7n���O�zn����m�b�����з�ժbͅ�-�ȼ��Џ_-0����\���NyHm�����U5��Lj�#�<�2brV�-�"�*�Y�:_��E��ς�xbO費ތ�-WW��?�:�nH�Q�4dֵ��_n���]e��A��O�8����r$��Zqs0�4����(f��b�%Y%�p�������x���b�$nw\.l�^�.?[�H�����T��le@�f���[��%7_�S��#�r��>�w�)�M͐A��jҬK<�t@N!�Tt��t����")�.��Z����>��Ł^%޻s��m����0r�%S˵*�;��\UQ��R��Lӂ��ٜS�]���<�nu��y�>�D���S��qq���fy��8Ჲ�U^E�U�Yg]��c�n�M�LJ��z�J�V!FH�)EI�G�����Y@��f��F���VO��U��0�m�̥��ϗ?#
H��D޳���&�^e#���MY��E�_\�<���a�mz/�p��q�Uo����/��A
"�ͬ�U.W���z��i�Y�_��E572t���x��	�$���"a�IeN/L�;�e[�'�����K�p���ܥBTP�j��77z�΁ݧ]���Ƈ9|1c�	��HHOR$A1~8�.�-�2KG���tz�V�"wb,^ϙ�i�CGγ�V�f� �����\�'Ib�>����}��=����%���q(�:pl��.)xQ6�v"/4�Bo�,\�9��T�WC��@�AEqkƆ~1[m�Jƪ?谕Hd���G~���EMM��	�x��L�&�ſ�dA3�mI��.�vrŤ79��un:ow-��>
��F�t&�u�=WX�[)��ie���a�B�=Fi�R<��[�2)ܮ��2հ���هw�>��-	�Z�/Ls��Ø�U���~���w@�e�
� /�?�ת���!��75U�������Sa�q��F�L��
�[�]�����;�?ɕu�ل��sJ�|[��m�$,^� \T����ӏ7�&ժVxQJ�>��[���\M�ՙ����d�إ ��ڴ�%�Y����o_&�smed���b�����q�8Y%~�ES�3'3���*p��LҨ ��Mޔ���p�0B�|굯;{b�N#
�`�{ w�-X½�p�ܜ���=�Q8���{�:���l&�h5~��A�d0��B���\QQ���a��\cp	�ȏ�l���9�6��� 	eae��o��ff�I����̓>�H��׾I3~E���nN�^#�Az�:�v�55�"٬�����������r>��Q��_�(E���)�� 2�q���0��O���4QyEI�vp�7��զ����bۻˏZ�Y��x��ЏT�1�MvC�UT��c )+�~A��� �����J]��_%e�W��:x[�]�>L��v��I����<ܪ�qm�AAjyPWq���}}X��>H�Y��켝�)���"I5�`_Y��x�s������3UT�笵`-zR��.���.:�: �I��9�b�}�8���x4߹�jg����I�g�����V�P���q~>#��J�c�{�B.Y�v�Qı�m
v�x˦���%D�r���� �\p��Cك����S��?�RL���O�-N��߻is	�=Ԣy���4�Ya�ۚ2�e|��d����L��z5�v�x�:�[�C��B���k����������yٰa���%�d���SR%�����^��B�re?�v6Z�m�;�Я]�)��KO����Y0���&�z&�.._�ӿ�O�������΃ �B�����I�K�_i"��,_�]�W�n�(�>�s E�r�5�H�\N�V�;2�2�-�F�b�)�<!���wK������4���t\����H��L=�+#��퍋�i��g��\	��)�ޖ�B���r�4��/�'��<"I��2�*!y��!���Y��� $hۡ��m����4��pd7.���c��F.�z�R�3��J�ӅI\
�]��`!`�r6�&Z��:�"�J�����Z ���7���I�3�52f������)��t���H��	m-�Aq� �af��}�>�@�
wk�5r,�0��/�1ʕb;����Z�?���)[�s	���^!
n��tzD���4�9q%ͯ��`" ���S*��w7�������w��'�r�u_��~� �#�>���nH��?��q�*�+�~M&�wl82M����?z.��w<�eQ�����(nf3�5�乸���x0��n:�iis3m�$&���C��·U��I�,��q+�ivK�~�1�[���|t��d���򂻱AG`��_vN�y5v���������Beb�ğ�O-�L\��pn�D�"�ލL����:��W��FvA*L�nGN������{�T$R���cXdX����H�~�@��ץ1��;K�tQ��?I���3}j��ۗ��Ű��Mװi"7� ��RY����Ͼl�7�R5�y�씛�â,�"���~p�J�p�'�f�Lz�R+-Zd<|��w�>�{�8`s�=NC�O�tJ+a�!�@L`=9ETC��̯��d�6Ö�C���{�y��ޟ����t�ńx2ϑb1�h����\��Ы\d>[0ph�h��DD[�v�v�4��ܷK��*���[�2�Q��	�zF]P^5�Jڋ�Ey$T<�N��Ͳp���*~<C��"VS�;zz7Z5�
����I�����>;q�}�퍨i?�_�-��?��Lw�������~>�G
��5Մ60\�v�=U����&�8.��vf:�#�&ޚ�ո�Iͯ���%��%��n�@�6���^�����M���;+j���`��ʔn�*���LE���m&��� }&���W�c2~7C�ם;�Ņ�2쐪ͻ/>.;����T	��4�B=�N$�ػ�_
�`{[�<�������}�gT��Ӵ�1�/˭!G��M5�8e6�kv3�xT�!�]��l����7A6�޵�C��I�6����0$�E����eE2+�a��?���6�h�f��S�фq3)��J[��l���E�[:4E�gC�f����� qY�"��_`77{"RV�9�v�Jz��/���f�x)��sh7f�/m�C�`�/�g��>a�����]g��)	�0�թT�-��§ P:KjNְkâ����"'Ϧٌ�Cww�����Z�;�̩m���*���U2�o"�?V��4⣝�q��'[�n(C��~ǭ�&�������6BM1Ѡ�鉉G-��!��6�Sʊ���Ԛ2ּ�Tv�@A�VO�c����jW�%Ī�Mu:��X߿sJA��nb ���E���(�3E4�< �l8��^�J7��;��_2i�(��9�r�IZ�5LUǥ�Ƽ��}��n�~[��M�p�`d+�l�/��ր������=L����_)���Jj]o�ٛ�$��8!�V���������r/^�����i���7/jP�_���������B�������?��ը�N<�>(+k��.����m��A����s�����e��E
|�o�q��2������ïG�q욳Z�+V6:���yh�6�}o��o�����Y�2�����I�
��B����I�#
&����7�|�o1~�q6�wjϚ4Ay������+�I�"*���f��ni�ȏ���+\SɎ�W���%��d�8#����<͒����u�B�m=$�<�V%�3�����)�����U����y�dĶ��iR�'�6��� �W/�'�D�M!�d}<����O������t~'�3�/w��3��L��u�m+���/`���Yƛ����_nYF
�� ��w�y�jl}� �!��4�#�>?{l!Tկ*�1�`�L��wa����S���̈�oa���(��>D=9:�XY�>:
�K]�=�7�ڇ��c���*�ttX�QL�G�&�0����M�����Q�Fs����W�\saRh�K�{:�ޮIS���iS6���hDEHWWgנ8�r���}B�I��:#�(�p1��4�[�`p�C���,<��*?�У-�&	((	�]9����ca�=�!(�54��}z��Xp�r ���٬���hWq�B;�[�735�ĕ�$��]��/�Z,��?��"�.֭����?�ė��U�c�]c����S\��,ׁ�K�¿a}��|���[;���E`G��������mR�M���2���ro����Um'Ĝ�@��j�K�ԾI	z>/��ܠ1�ۃ�:�;����d\��j����<!6J��T���h�KP]�`ߗ�Z)���Im�a�;�ۓ�������3���\�iV��Z��n2Z�ݮ�_�X#���PAN��ggo��7ĬB�#1Eا
l�o�v�/�ؑ������`�C�Xς�f��B�L�r`z����Y����Z�K�m�D�V^M�Y\^fz�y�����b>�u~N� Ұ.��|A�����(�]�b9� �G�;l:媳Gp���=�B�j��oN��G�!�:v��i��?1j�z�<���ì�{�y*T1J�5����9O���>UUԉ��ׁ2������QsЕ�9�\{��V5���Οz�{&�ʹF�9�Yp�ٯp�ݍ��;�3�T���`@&g����BI���B���1Z������V
h���vMa�������
K��{g歜��ֱ
��K~�����y�7_%\���8E��5f�2����B�Ҍ!����"�Q��E����2$-ݎ-���Ǖ���EIU���~�&kQ���V��e�Y|!M_������֪��Jx����d�T�}?�	�A��c���=�րc �����'�t[���%l�ݙI��P�,�U��#�<jT׸D�I���p��'Ox��L��u������_��u�}�n�WdISzKU���G��K�v7�ʐt��P67؀rE�����>%���L<��wMy��1������+��('08�V+Y�(�3!/�~$��AJ{�d�q[�����ע\�M�	�^R�p�Zӫ[b����BG[	�stP}�ܹ�<�ɇ覄��5��P9[��*�����O�I�q�N� mFWO��M�)N����W��|������_w�L�Id�|��]@�h��_I��Kn�����9���nJD_�qC�?������-�n�����ߏ_v?!rX��V�GQ����4y�O���O�����p2���;r�����`UX�6v�q�]Jʄ�S��'���(U��1�hy��>���Q'���6�q (E��z�����&Fsb���c�<�H�K�M��^%�r�VNq�h�p�wS1u�>�2��׳��_�����08��(v��H(y)�G�l�����D�S���o����wYY꧊:�7�G�H$��<_AyZ P0aFy#�+��@%0Y��ٹY��U=����c��<�b'xJf��St�{�s�-7q��<T��[��׃.�L?���I�b��=%��m���ͫ�Hb E:W�93���:�O}¸�V{��˃��p��j�8Y����Wd�R��^+*��8Dr�/�,Î3I�&��� ��uP�L��0�q�,/��ai��i���z�&�xq���J2�Y������bM�1��AoIH�!8#eg��=ջ���0���QCtI���~ƜuыRC���t�(�v^g>�)�)��AB�Y{9ŷ�7��loW��U��ѱNw�
�n��-������ɑXٍ���S+�<Y`5L����\�՛���l���MRI{����A��9��e��WC����)/a���Q������!�>�3)Z��?�����`<����>������S�lvύ�����э�T��,eL@pV�K^����}��2W-=j���U���1���^���y���>1�s^ְ�׊��7L�w�ldrb���%�H�H5����w�%m�Ն��)}f��	���X����G��X�؊e?㾽*�=���:��]j�����p{A�suu���x�>��ۘƾ�q0�`���TDet\>�)��H�0�͸���~�/�y~eK��Z����v��3�;�L5b ��{ܻ�v��'���,��C#I硊����^�����f)����ĺ�{�7��f7���'�Z��W78��e�9Q��Q)u �Y��ʱ���DN��*dda��(�X(�a��j��J�K2��kF�;�J_�v)�s	g��Tx\�i��X�*R%���T\a���k��@��L�P9 ĦePrѼ����$�����K��q�#�`𔛜.�I)�/JP+��P[�(*/���b��A�We�w��[G������͊'�o�)B��?�`�ꄓN�{x/���c��G�[�5������'�&*���~�<SRI��F,E�{������g���hK=j��T��C���frWxl�lQ���אk�[�al�D����^?������nݰ鑤ÆǷt(oq�-�ġ]�?
�� ��Q�y�j~E���������h��^��ty��~��;���Tk:�W8)5�9����|��`�fo��b�����Ew��l[� �ɥ��tY�th�b�y��j���L�Ҏ�>ܩ�)��=���ła�ȪY��hK��3�t�rY{ҞM�f����Eeօ�N}y>`��Y��7�@O,#����ơ&�~�z��)�bE-������^nnn������-'o)����;��-GCh��[V�U�I�=�z'�R�������c(�>�B�	l]��<�~lb��+�\퀑�9&)�~�F8W[�rԟ�Jh�E���|�s*��~ ���W����3���O��5�vX��.s�.[^��n\������~��f���b=�|;o:
��ݬ�2ػ~/�P�%�)���B4�t_kQ�xU�UN�tI��ȫQ��ݳ��nA��伽��[[���g�u��B��^g��r�I��Eɟ�?FG�(S�h�9]hc i�K�WFu�M������	x4�vuR��J�59ץU=|�@� 4����j�	ĝ��5�,�AH2Q�̠ix��Y� �3Z��^Ր�V^-�[�CZ�F£��Ͱ���G��۲%`xx��E�0��%g����^���,ag�� EZ���S�� jGX�<v>-*_��/ǉ���*�0"�B�\�>}�O���f�7Y��2@[����Ș֒������7Q#}��K�n���gn��BAVy��oO��g����Y\�������ܬO������Qg�9^�1��B��??Ce�ʝ����ʾڊ��]
���PB��S}vL�hR�Jy�@�n\� 
Ʌ��?9�.�v41#ic^�<��h<�B�D5,�_Wy-��������9��Q��az�l��ǲ�����(��nf��I�kiJ�# ���A��3��h|�cnW��P������i4T\';��Q�O��N�H�1����Уv��H�`�u���;7����]��,<\\� q��^H|M�.c�9���U�N(	w)�#��g�����v�LJtQ՚�|���3��ӛ����ŷ'���3�����Z�#�cd�`%rd{���粄 B�	�T�^>]�;�ˁ5-�G�{�o~5���n2�Z�Z)�`k��҉�?,�j�ݑ�5B�/\��ڟ�Ώe(�q�偺 �@��#���_����1�$��	����`���;���ǡن�@0�oy�c<�J��y���B#f��[G��O_�Ub�j�ه*��G/�ٮ��߻�3��~O��Z?n����Q8� �H�c����Ͻ��|�,�o�iJ��sWq��c���g��,#�}�Z��ﻹOR�/�z�UO�ܚ��Q� ��a{D�� ��\=���q尰V9�sƍ���HmOi���w>0	� ���5~�AƸ��B�*8#�0��VJ`RJ��*���^�iH�qo�3[���
{ ���)����q����s���`6�����AA�� s��#��q ş��IQ��CH������F�>]ȷɕ����Ћ�
�����^��ޞ!�ª���	\1K�^U�˝t4_��2E��nl$�bo/zз'uA�Q����Z�׏�fm��@z-���G�YFE�Em�e�F:�q@@���;��n������[IJ���Q��?�%-)��������v�:�޽����=gQ`��/z�C(wuUR(�"2N^.Wͦ�D`��h1��'�Z�a �R����'�-�QD|v����w�=�}�&4ϛ��(�vʇ�Y�Zp�\�ٽi��I6�~�Xlȵ%}�eiW4���߿��[S��/d��<�ȟ�'�J�	N�z��H��sR������8F�Fђ�S�N����/Y��k���e}/�4����(<���y�w��&L��#!!����&�g]�����k��?�7_���	y��{g�����Y0םfu]G�ʡ���g�r����+��o���@n��~o�ç�w�hg�5��/�sR�A.�}5�?M����~�w�ED��֜�a�C���K�ҽ���q{3�D�s��A���j4fq�_A]P-ks�s�<���#�i��������������WA���gw6,<Rj�o���Y�5f�wyc��~1@G8�v�w�N����h���_���\��ȌU��S�}Z��w_q;Q��J��W/��_��dv�	�w{'"���Y@�?,8���i�)����Q���A�@��_�ǗIw����e�'ޚ��KJ(��g80�һ�J$�F.+�Җ��!t�{ ���T�dŪ�'H�9�3�3�]��u�����~HZ�<�]ZY(�=��Qe�S���K�����`Ք^�r��q�����8Tˌ_eg��r�R,��cs��Ȑ�d�ͦ�����,)�i`a��Ѹ��8s�n�%�"!C�ŵW�X����#Y�qO̯�m��
Or(�;N��Xhvz��c6��G�>Y����Z�+*D�|i�b��u��)�8��Pw��nmo���j��e�V�犸X�,���C[���=\�vȍ��s��n>�5=U���O���~Ǩ��.n�K�OܺH�4l�R'�0���X&�+y���V������ձ�gԻ.� �{j����2�T�-|�%u@�i�<3�`=W��2k�d�X�Z������Wߖ7-Զ�iE���1m��t����܄��k���s�)�\
���]�4#�s9:�q9YЫWSed����"4	g����4^��#)?@����Jצ8��%�V��=����^Ԑ��Zx`�<L�,���=Q?p��KPZGG�*H)3e���(�l��H/I��b�>_o~�^�}��t��&���锝"��+�"%g��%�*�%��VL���S��+��>8f�+��TcCǐ�F��T�y�2���_��v��/��e�Q�E�/��ǟ������? w���?�m1�uXz	�it+�j'�2����˻��b�W��E��gŻ��h
QҾ����'���%?B�_�"�6t���P��jZܗ���j,��=JK���/���w����^���-e��wp0_��a��Ct,KL9+��'���jw����ʂj!.��67�`h�f��f���{$��)YV.d�D�Ň��]�n^�!
l���/�� *���"!-m'Sⲿ�5H��tm�>B|w?���1'�픖����
 <�,�`��~�/���c�TQ�F�$q�}7����t��F&VAlgǾ�V� I�4Ӛ����j��(X��m5'���vI4�?��@��.��Vު;x�� _M���;Q��$�m��Tb��K�?~��B���[�y��ڀ���
ad�ʳ,¿�%>���'�+
x�s�G$��`�>Bn�S�?
2������I�p��{yO���tyy�x��U ��q1{��LMm�� M�mdN��%���Kv���2�86rTC,x��~���%FQ��t��ؔksً7���Mr ����]���0QMTh�������%�ş�[1�D����)?�u[�3K��Ͻ�x��Y̙Tj��X���7���P�[x����(U�Oo��z�	���u�f��^�}n��tC¦�x�e,^���\�5	�����Zd�C��Z�F�56%K����e�/�2#¸<����e$�p��9�gRxK$�<�mhh��	��]/$�q�6���ж8�����J���BT�*�hf�-��/<���(�{����D���h/_�\�r��S����H`	�9Z4�A����՛��� ��I�>'��=P�W8�h\���^�o�?�XC$��]E��DGK��|ǛL�͋���H4~0T�%C�,��A�� 齂���~l�'��K��ϵ'�J'+ZKѰD�����=�������ѵ�	��Os�D�|(�
����T�2�����h����й�}�sE��>G-��L�l��g�	�dee�	�k]� E��R��
J�Q�R	߰��t�Q�5��Ih��Y�3��=�d�_}5=[Go��$p��Dn�Ȟ��IS�!mz��ސ�<�u���J�j֩4�8qF �{�|*�� ��6]�-�����}��ۅ�֟�^��袤��E�e�;v��Ky�{��ӗ��%�n0���gþY��\R|e���o*˃��NA��U�$�5�f5Q�������L3>��3�b�痻;}�*���i����PNd�o@@ ҿs���3��1�zl��O�U.�S6&қ�7By玟G��+��ԟXE%�A	&�W����14^���y����nվV���.�1�&�_�M��2>�*4-��>A½,q�Fx�(j)�(V�?�W��ۘa�;Y��"t&��{;/E��Hl�'����8��zڋ|��[Ɯ��ut� G#��}�M}p7j��ٳ3u�x��;嵳�th����9N_Of�J��O���,^��P�o���b施�Q̜��u����"l��B���t��{�؂�y�.쉜�6E���Zs>��+p<2��50�sY)s�)'��"��_�[sp1�M�͊$IP�M5y��)��:���
��L�>���b��>�k�S,1��𪭭�Ɲ�gy�w�{��/�������A�C��=A�Y��J3���8\�7VW��������A�H"G�l>�}��Xst��/R:�|D,�U��)��; ��ٵ�4 YZ�>\A��0(�(Y��9���:jd8��PA�I�A!>
� �+o�X����M��I�MI))�d�i��@��0$��r����.[w��wC��]G垶�gV8>1nMT�i� 2Br�S�Q���Fߥ�lPﰬ6E@�e�kvB���-��M���؍4�k���}s|a>�Љ���9�4%b�q.���2Ȃ�o�A?C8������m��),�y<�/���s�4��Œ�C������ڏ�+�X@�,8OR>b7dcz���qmG���fHt������<����t�4b�L)�
AL9q��i�!��9`ݼ��Qz$���
� @ '|B��S��ܯ�z���'6Y�X|����
�y���@�����Z:/B�;���"�"��!"�Bɚq�s_K{C--2喇��f�tLc��N1�����c-?�%y�����}F߹Ȍn&|m�k0�R00���S���c�Pt�3X��>�Dq�P�"��/BmFq�|!`d���)ذ�	bV�49�|=i<�Dv%Q\!c� ���X�$��i�&ПY��N��m�}��SQ;���Z�X�!�эr@��2�C%0�C؏5B>eJ�&o���F�Z�D�wգ����E1-*���)��n9�|.�w�S9��������ZB8֮�A#w���BU��c"!'�`'dLT� J�/Le���I���{�m���Q�Y&�K; z��}gNQa�����먩~Û�6R��u�!�Sv�tt�Y8���_�Y�lk�� b��T*Ƚ�����B�O�ϮS�l�����[X��\\�r�s	h�HHK��\���W��OXu����,�f�d�����A[���8=�N�V�g�j����n�2W��c�o_VJ�"�ww	�2������88 �7	��j��_>��e�������K������^>���Rj\�����oı\���{�o���{0B3`�b�i��i��Wb��Zz���\-S���]�VcB�r��Ƈ�#�ӂ{i�KE�y�;!s�04�quI�c��o%?x��#t$!�]^*���a�����K�4l�B
�>ƈ)�2*	s�/�}Z�8�x�ƞ#%���G|�1���"`A�eSw����$�2]�������u�����<��b�*fX'��W}?h$Ip����An�Q=�b3h�� �/����@n��.9"�Lt�a�=�՗E�Ab��	�eU#� �8�gba�S���B�_51].��Z�ǡ�vĹ�˗�#=۞�vtϚ��'$��D�����HR�Y.k��uO��h��|�p{��:��d�u�RE\�a��]e|4E�ܪg��BR��hb{r�Ŭ_���#U�x7�{��@�'Q_-�����J��_�}>��!Zz,�^_��IT[;��a9�C"��y�ۭ;���|Ā�P!��t_�K=��L��d}�4n;������l����6�٭oA���Zŀ��Њ���该�y��xw�2y���{k��I�?�5�?B��a�ާ�dDV�{M�z�$���撨X�{�^]�w����dz.8�X���� ��()����~��q�J'���`�_��h���iz/t�$;qK����ޗ ����M�����\�I�z��-;�/}>'�������eNX/V��I]��}$���$Δ�M��0�MQ�54�[��^�n�4ɐ��`���P�&�V���;7�i2��**MOn�(����3��=^C9�yp�����C�Q6�����t7�
�^���t7PV�K�$`�]�#\;X�(�����V�����:J�˲�s��gLK9 \�
$����
�7�rJ3nf
�o����qbh�m�eeQr{Z0ź3��=Յ�E��E��R�%_^4��:H�|�ת�U�����aP�]�I'�4.�wƛ7`/�<jx��ڏ�A�4\qG�5���hq�6:�^)T���(s4$Lׂ���{�������U��o8r�.r�u��7�ם�h����c)Wu<��?1��Ŝ|Pt�4/60nU|��/���oQ�$1p��lC1�;IlH(���<
:O$�8
I>��JX�M�gǱ������fsasa9z��A&��:Y<xEn�H�v�8�']ܞɸ%�
��E�ż1�Ϥ�y�ܛ��MA�c���*&�?iў�)�k�(�)�oHݜ�
?K���_���7UF�����I[����N�%���,�Șj>���{z\�ӏ���ы<�yU����i�_#6r0�&�!=�`����{��C�9uDud׵�vQ���H���P0z�|b�ᤡ���}���n�<�:R<�� �hz�x"~�A�%s�w7{O�ҕ��J���$�db4�C�N�7��A��Ʃ���(���I;<��ʼ��nڇw�}-�Ƃ�Ss�����:�5�\e�ᏻ�I^�յ�@���T�~��z��Q��uhG��{��K:�kT�<�2(
�i�ﯞr�]��0��ݺq~t���cԿ��f?bv�žXX.P�9l�fE�*>)4>7��
Uc�Y��(��l��|3Tr;��>hؿ�@�92)�A�.x���(;�C	�T��-#��U����w/ċR�3g��
�j���+���G/��ֿ�|��(5�:��ɪ���E�����U�$��v�i��ͽO��QOߨ)�%�xU����|sz��'�����o�K������{^r�����X@���w��ck�=����˥��yV�cC��G��[	�w
������CҹH�;�w*�v5�������5����r���JϏ�FِA����w<Ї��]��\�FW޽�k�?1�DLSh$��-=8�1���߉{XF	�G�!�	a>�v�4��c�d��aI��1^�3��j�[��7QG�=S��8��8e���W)T�]r�}|�zt>?I�M=�d�2H����3���w)�֣��^�v�E%��*#�eFi	�'vΊC�5�=s)�r���.��`�ɝ��ɀ��`J1�a�!@=�ɴ�X=cLXőf��
�+Nb�A�����j>��]��Q��K�똜��x9����{����S��=WG�>�o�w��魔3A��*�kݶ�@���h�L�15�R�s�(�����FV%k�/��+�F����ܨ������"�;;�Ԓ �8Ҧ���!B:&��6V"� ��,*~�|��`_�u ���c{��>:�s��~]�]v�46B��4Z���{���G����l�T�0����T��t�>_+߮:����?G'1��ͽ���l�dT���q����	�D�e�d���Nj��·כ�-xl�-)q2,C�鴐�^�����"I���n۱]{�h�t\Q��q߬��������x���wY����z���L�hb�:�HY����x~|����p�.@,��>�`������L����*{	J���ԡ�����ƺ�)hʗ���\y�<g�f�H����p�S�}�;t{���3`Oa��[����+��?��]�p{�6i9��uZ��8�؍κ�	6���t��!8c�S�k����iy#dZ!�����=T�͍��h*h�9Li�Z������ҋ�h68u]R@���xbq�i�y0T�[�ݲ��ϗ���x�`]>3�<4Ά��5���F-dcn� ��[��Q��u)h�=���{M�wV��4��^F	,U�����z%��/t�<�#ɂA�k��Ho�A.(��ҧ�N<q��h�ئtD?�_�w͉oQ��qh�B(^�W_q܁��C�k�=UD��)�v:S�:��.��5ե��|O4�/��Y�� mt�6>��!�@�D��LF�t�S�>�5��q�C~�^Y��k
X��������	b0��P[n5��=(M�jsq�:��5p��:��r�g[�Dk�ڭ����!"�"-ab��b��ht�Й����86�"73��^@w-{���'����n,��.Z��?�7���{��]K3�){_G\X����&O�z�'�j�e�u@B�;�LmlY��s]��FN"�{7�gD_��|È|v�L��ӟ�*⏠�ȟz׌���������#���pF�&l����TQMq���	/%��$�~.��z���G:����5ȥ��0~}.j�v8\�o-��7��7G�ߝ1�"F�z*�r�8;�c�
+��6���D�,��t�֚�|�U �|�KZ��#��vXT�Cy�I��j��Y�)���*���8b������2r��1�=�ӥ��ܤ��T}�Y���'c��y0�uB��O[���\�$�Цl3�F�����fnrW߅���n8S�!X-s��jWJ��	j7���0��$�� �KO*k�!5���������z�
���n�����G�Q.��a:�߰:H��r�C�A`N���j��X2#ƶ#R�HÞڃ�-i�R`D\n���,U��ڕӽLQ)���Y'�z"�m�5�&���xL�њش������=b�)C͎�;�Ax���>�.�A��Djgy�{";~z����q��ˢ��uhA�Q]�O�I��ױ]B̅2�v7��SJ�z��j�s�R0H?��h���'Uk���35�~��<�©:rO
�X���W|�f��ݗ=�4�K���la��'�<�o�ڏ�r����gO8�� )q:�O�;;!{�qC�>XD	m_Z��n�:>�KYW�قf�:B�"��*�42�m!jt��O_�����v���Y�[>D}��4�;��Uz��4�����a�C�GVG%��S�������a�]�6H�"6Pβ�Z� y�(c�)GA�[3�
��F���?| ��m�
��L�Ơ��w��������?�����B#Ȟ�H8�,��F�n��3*�C��f�=n�n/%���懳�W����$�?���9a��VU6~��4h�n����=y\F�č67�MbT��ݻm;���JRֿp߾亃��9`%�@���1�	+��DQ�k���s6�@[m�<k7��d�����d�οZ�,��T��;�X��qp�$J�uF)�D>qY��̗�\���ן���R��魆���Z��5W���kSBЯ�b�$��[�%�.��j�n�>��/Q�Ά,g��SHa|s�1�V�5B��a�b3�9O�:��;��p��u^��ػ��(і���Kpv�Ix4�n_���*��Eᔽ��@�ư����L��v!<
�)٬�߳��FȖ�B��(�մ��R9LJT+�l����d�|�d�(�b:؜��q�v����A�g8.�.�ڋ3�\���4�v~����E�ŗ��EVmr�E?�[=$�G������S����(~�^��Ku7��$�J#����<.��7�$}�U��J�&��;eSEd��x����[�>����셎������ќ	�5�}�!�;�vُ���<|� ��]_�p}���<��ݿ��)ܔ�*�����Gjk&GX	��)�p�2�>����a�֣���l��(^Rם=>Ѫ%sE�&���w|�e^��E�ӹ�
F�:��@��~�g6�n8
Ïe�;�h ��>I-�W�غ����d#Et��^��i`2�lh��v����R��I��������
rr�R�&�_t���mC����hx�]8|r?=s�=v )�l
�y�k��D_�m�[�c�i��D5=A�rTD !-�e�p8��䂹�,�p�ش�M���g��q�X"<�C������VD�������j�
:Tz��e�X .�!�(���Fy�F���<�ҔE���4�zv�<�jLe{��ŵOy�cX7�n�g�KO��/%3����m5ӛ���~|�7��YVC�]�d��ǨP�y�p��N�]�沝[�"�b�Ǩ��$3��(ꍞ���5� ��y2�&������f��"���Pz�ƅ��x�8�i��|��nG1<�#}��'j_�'n����w*��7����8�ʆ�gj�ϋ��+��*�c`�^�8HIHP�T��s{3�m>���"�+ݢ��'s@2;�B6}m�t-����v ~]�F�EV��B���S2^�����E�����[�ߗ�U���7�H\`>Œu�&��` ��� :�T�}$���
��<Ԍ�!�[_���V��=����|� -���0P#D�4��7�
B'�#�;1S��=�����f��Ekr�i��S�%H����3�&�����5Cl8��@��ד�����+����|��lZ�q�]�����v|A�]>�Pd���c�勒��YӮE�FH��n���|:��:4U�ҽ]��o��#�裝��&��A�9�?� -�g@H��)_�jƶ�mDx�v�d%�\/���&�7�SR���o0�%���q��XN��hD�v�{v���pV�|�8�5A�l�E�$Ǔ�1���o>�-��3�n��F��SUQ�	�y����
48W1�5��-��~q�R�>�4M��|P�[p3L�	 Bs'�W�dx���.t�7�y�}�i�򴷧����అ�ؚ�'+Y�4Ij�qm�R\6yL�m�$�=S�d�_�wp�s�>�v��}���|"���dCǾ���A�� �(=����t���f�t�Ú��ț��ܕ� ː�����')����?�g۵W{~��tO�<%�e��9?�T�_�5�=A|�j�n�X�[{��d��휔ٚ㮙��o��,�o��M��j���L�&��/V>+�M�"��V�����&�8�������Rٻ�]���⁷�wmXG��m�go������
m'F��'����|_v4�pA�m;��������xԀ =��dI*�o�Z��5��FPÖ8�ૠb��j���

ݟ���a�1�R	YY���&���0{*|Y/�:���|<3������w֏�s2�W:�P�H'�[�n\���Ӆ�^���ڂD~���e.���$��}�ėT�`�j�L��}����r�{��`��R�_f���<*>��'�yb�6Rıy�ץ���Ѩ��b��^p{�w'�3��X�R��@��jE^=������:z6�78��@���
�E�JՕ�_�����;�"y�h�>,"8�O�S��i�A����R�E�|�i��I�<N��16�ͦ�<:��S���Z�Rh�[���'���k#:<84���!s��K���s:��SE�Ǭ��i�����D�� ��!��(U}���4mҠ�i��B~��3�ͦe� >#M���$k<��v�<���XW���&a�;7Г��y�����-Sα.t�A�������ק��*Y���o���������,&D�P��#�4����1�D�p�T����](��m�BT��i�P�U)g��z����ו3E���-W����a5�w��@�)V�'f�@��B��2�ɳRO�`C���T�06�*���) �OS.dk,IP��a�rFAs�����T���U����Ŀ	îy���l��)�ؘ����~8w>���JO�-
Nq�G���n�d�r�
�J�oj��r�J�~����p3
U���Ңʔ"������@q�V=W�x���1���e�Az�#����f��.�]md�h��H��/f3�����ٵƣ>�"�ʴΏ�r�H�
L9��5s����N���p��R�����=��V7�2�Э>��.���ّ&�pY�B<:�����uYl�>ft��x�1ɣ�DPU9�B�O]�Y�#o�8��3D��'�t�:[m)������*[�� 
&��B/���Y�SJ���ô`���)O�LJkkm�L�;��'4�eP�@X��"t���F��%n�P��!5�u+)�� ߆<��0��D�L:� z<�9��	J�|}a���â����Y��O���d�<���*˱��g,nA�&0F�v�_#�A�&�=V���o�1b�6�婆k��T��R��:v=��x���;�H�%<\�J���?�яo��	�66C��E{B�����RW��#���Sԥ��ʦGXн�Uo�M�l�~�=Q�=z��>�w58��������_�É��u�@T�O<O��m�t�8E�(��}*�I�Ӝ:�j�\y2O//!:P�{YA�/����J�~���v���n�K�G�~3��)1�b'�Gud�Ѷ+���ԗ�^k2mn����6�E���~��P~��#��@�YI� �,��E����}�����m�|�x�5���$%bi������0��M6@������8�ę� �K�p��+)��� �FK,���$ n��S��c���%.�c�&�ф��4%�Z��f3�D@��3/����gIs?�$�OlkV�AF�4�5���9�����E�_O�2�v؊�V�g'~�H"��ي�\��\�GVΫ�����LN�]�_j��F�Y���ٛ���-#&��TE���x���C�����I��uX������@N�025�Sm���%ćh�h<��x_����Lk'���L*,�v_4���,72�c���X���r������c�1|��.���A%�M92�^����,.˅���i�����X��
w�^pƽ�*�)��3��{��Y�L�f����3]	�8����B ջ#F"���b	��/�{���o��9�^��L	<���4�^}�ݫP�s�|A�%0��UKW҃K�4�Yth���[�(���7��K�YJr�#��lP;#dl<*
����ӟ��~�}uIss�'��5��1n���Cϩ���6<mx���?r�dԽ�j�ɻ,��,���GaJ��ss˓����m�>��=� �7�����4-�����$���i~75���wr�th��o��.	f�$���d2�IyK����]�>|��ˍ.^�Q/C�S�$�|j�:��pS<Ÿ
U��o��Գ�rA��+���tB��s���__�Z�9D*؛�4���Y��D��\�(�M��S�=o)����a��{�����LW��Nd�fm\-\��v6���[\�-��ǁQ����E�!�^�����x�	�"E�����?[���qHu�p_��T��.�գmv���x��H:�:�d%�ǟ�`�A�eo�����W+�p?��xFIW�|՘P���HU�~��y*�����#X�$X�P)q*ڲO�q<�<TG/�&��
��F�G�g���A��AF��^�߿�D���0�.;׿�λ́�8�kk���_&�c׬����Kw�L�L��v�����Rt��ѳ�3k���_���62q6E����K 'a}�G\�xJ��+�{4�r�5�Pd��jᏩJY�9�Rxشm5��{i��]X�W�7�շ{stG�SD�^�Q+ɛN�O�cوƧq�+8v���)���@b�����AL�Q#����[��#R��ׁ2L�V�7�8A*DPZ ����+���-s����#lP�t�a�ium��cj��j0sa�����7�nE���3B�	,����3#��[���ط��1��x.D����=���׎	���h��x��l�:��'qL"��Yb?�k�kp���a�RҐ��\�G�@�b�P�� ;OJ!_,����z�"�.��8�Ք=�{��}��5�;�����(�*~^G�e�X�����!�u0�m�&�T/��: =�C^�*#������-ZZ[[{%ķ�ºȒ�L���^�B%���R;\�eZ���9J�����zc�.�Sk������2Z���}�Ͱ)։��N&�
rhZZ�k�p���9�Zä�B�ن`Qh�;׳v&��Pb(4�p_��^�E��I=��'͑�;�]-N8��@�C�\��`��F�����i�;t����S�e]��:Ϧ�t=�?h
+J\ҥq�Cc^zX�h)N���)�1� 2Oݎn#�UDY�y�}�L&�sc��`S
��g��#�h������%; [�d1�\�c�p����U⡿���N||օ���Z�;���3�c�DX��s�����T卺z��*=�h��~�9�{��_�Qd�pX��g_L,��M�B��z�M�P��9L+nf�pZ��w"�A�K��Y��§�bW+1��/�3%��k�ꡆ>@�I�Ϫ!�oVe[�s������ڋT���K�g<[���m�&��k��s��+���e���l�9jZr#c!8�����ףcע�,�Bx2Ѣv�<�{���:1R)��b���:5�/ ���΀�N��D��}��v�R8'����j�y)�+L'_��}���1�1�ׄ��?�� `_�u0���0�c���������>�8	�9cz_RRy���^m���A�7d#��
�]����v���[��Y����H!��j%�r!2��\nt@�ˎ���EJ�t�w�2��� �����Bő�[�	��+3\7������顱���_$��Q�{
���K��n��K~1�4����^ڨ��wb.�k�Ţ��]�䶣�L��#~��U�-ut�;i�m-�������8����Q�ԗ���E
������G���=�U������{�K��X�.�����o�˻{��E�4O�r'k�!��H�c�7��FYF`�+�?��1u�U��GɁ;9�?��[�<r����;�l�I��3�#�;�鈾	�]C_l(�x���r?�y�ԅ�uK'w�p��; >f+�	O ���Q>��z9Z���a��<� �Nj��7P��%��)��$�p)������>�&�7u�w�h�#0��S�B˿i��Uj���6r�JJ�-;7Q8���c89�]�*��_��Ex�7Ǹ�+o`�p��1ĢF�sZq���oP% �a��G��#o볋m�ne4�.ME��V���Be�(F��c��K�P[�yH&��	�����Rɔ*��Վ�ן>��~�0�&��'���>�
(�!����2�,�e��1�C��-�V�V[�ٚ����.Á��Ɔ��M$�C�K&���#Zz%�N^��<���/U��]��}q1\"n�m���w1Fk߰DY��,ʞ���la7@�oi�zA`n�,�V,�RA����{/�p�U���LE�����$����(ua���sOiR�u'F~�00�9���La�O�%7�d�H�!f�7��?&�]Jar��HF�#;QW��f-p��Y`�;����;@������-�'�NUN�Cպ�E$�,̥�|70�2��8��z���p��K����6���*<q�fu�_,8�[`��Ň�ތ��w{�V+�ȼ�q�9?����'Ǎ��2h/o�hQ5�`���
;��7tx�X�L�;���0�R���*��7;##�
`l?X�Jݲٍ(W+�D�m���C
�OSh�2j���W��{?l�:�{��8*�i���)�?t�I��Utz���s�DEE��c�����e���8Z(,��R�x����3V`9�_��L���z5����AM��,�WM0�[�Q$�
R�l{��HDkLK��� ����ؙZ���g��D�s�4��>�c�Ƨ���x��_8��s9�����¡��
��0	���/�sub�6�I3�z,!�yb��u�N?pE�S��7x��ѳ<�e<D{�$�=J?�[`��ǝ��qݍQTXҠ�7ƚ�H�p9�!�K���І�z�bP���-�qCRv����Y�~���a����efR\��Ce�70�V7�T�nԄ#ddȯ�$Йɽ�r.�/�;^;ݻ����G�\����7@d�������./u��ќj<�����/�58�.���O�:�$ı�@�S�oR)}���l��!�;�FR
������Ҿ*�-�%İ�.�7��)����A�>��N�� �+���rP�rf32�x�T�P� #=Gv�dY9�v��A/���W���J	��z\���G��Y�ϲ7�4:����mq}��@m��X�?����#a�?��7G9`��
�S����^�DSmV�웃��4㶩��h/�����d�e��c6qG-�W���*�{3J�G?8�>���� K��u�5��ʁZ��?��զQ﷿f�`)�V��}f�qc^!>r���H���F���HC���g�g�"\�;!�S���W�ϩ��.��qo���I���Y�{�M�!/Gဆu[s��FM�8�s�v�}�i��1�c��"L����1��d���<�G� ��Won�LI��6n���7�ȉ2Sf-^
3�y%ڙ �'.Wn����x\���_6��]�W�+ܐ��}���몖�
Px���_��X�:�(��'޻!�_�~KX���k'�M"��!�.���@����e��4���x���Wx|H������R>� YB��co{���E&;��k��G e����M~�P���K]L"kVVmƘ�"7��釳���	"Izu(��C���xrSaB3��]�ΩsԿn��s�{���� ��D�!�ž�!�Z�� �+���<VxA�Y�K���d޽�"�',W�g^���?��iQ��!/�ɿS�-7�3 $�\d���/��2L�KU��qr3���s��KIoe��|*0��X:��Ϧt�ؓ<	�f}z�v�!m�%��>FeZX~���@�j����|�'چ��8�i�����S_
?��`:I����f��m��K���׹N��DV�4��p$	��7;M�dT����R���o��.eʵ��D�5j�G�.c;��)A<*/D����g�Ici��(����Dׂ��[��>��7̇���(�1�?z���W;C�sDD���,��x��$]��:M凱�V�7.B����������K��fr��&��n�!n���i���`�&���*-[r��6�	GA;�.�j@��Z�J�!�D�p(uP����(>R�i�m�Z��J�X�Z�����}%�����gg���:�J؉Qt��ExJ�Li���������2L�K�7h�8_�㖚�`ԅ��ȽB���H��=9��Ie�"c=!��r��y�ˏ?fE����j�I���/s|�AgX|<�H[p#�p`�[��㬱��L<�����A��?�OjNA	6tWY:���@-&?��پ3�X�'sA��$�4h
�I0��H��5����m���d2HaE�ozRǑ��K9��ْ�B
�_ 0�~�@&�m��e�^WO�
�E�~B�R��s"!Y��E����P��XY*"ty����nÔ�����IC4 6_O����_E��ά�1�xNNU��O���q��|!1W���Z��c,oh�;��p�������9�!(����*�XT΅��R�ҡ�}/*6��n��-G%�}���E*�a,j=�ϓD �㼱��y�I���2�>��F�WV��s�`q\�|F��J�u&�,������k��>���%�1z
"�%���)�hāG)  5��QN�tHw��~�����k�{�u]����D�����������ԚKf���0}�S^��DE�#��C�Pw�-C-�������
��4�����"��r3I�{�=�.JM����	~Ϛ��έ}�����|�5ë�(��.���{G����j+��'Q��vu;�BNK!SN�gn[���civ�����\���Y�7�5�z��� ��	��X@pY!/�c��8�uh4ѭ:��}w@YyboBaDX�\�o��������[G��2������
�s0�T`m�s�> 0�z>�?�5�5|
����8T&U�H��P)�Q��p~mI�,Y�V"�\��_�g�]��κ�M��J��&�*�����M_A�GG�+ˬ�� Y�i�жP��@�\2.���V� �B��jw��y-��~O�(Y����|󕁁/��_t%��/>�V��|`��8SI؂���)��"F$���=�[��1d���:(��%j��x�3@��`ֹÌ��t�Aظ=u1�(��*^�8�����}��!.�2����88�i�"�A���&�6J��N���=;#�������t��sx`k��ݺՈ���WO*��W@@�^ �Ōu�D��|���u]_%kU�&π�o:��
�%i
ڥ���-��iȋ����+��WEE`��\j�C�*ͪ���B��+��띲��o����O7�v�C/,Tz0c�)�l_��;�ӊu�T��k��0c��M����>��0��4
��[˗ʢ*�AAaj��l�ITܖv���[��%��JP2H�D�.)E �D�m�ap���B�s�*mb�g,	��;��n��� q�폱�Y)Ӈm��z�+�\��340��ؗ ���c6���X�J�������������x���>�j��|�C(~�Է�uB?�cG�����٬{`�� ��C�� ��4y���^BM�K�gYU@��҈��Lo�]qq?�FMG9�\�k�!A�EOr�E"�!d}3Ez�{J�`�l$^ ��N��ҥ -}�W=`��~z;�W�s����Q��3Я�s�����ȿn*��(����V7*���XoĊ�I���Ӷբr�x��Y��(��H��C���C�r��]!�5Jm7Ϊ$�ɛx�G]���5�V@B����������U$T���: �Y�S�����7C�I=�k?N谬_�d7|��f*F�C�E�|�F�^k�2� ��F\t�\v�lx�7@6m�[��c"�uXn�dmJ��1(��Rӑ߷���`,��|�Nt|ɪ����f\�hQ@4���m,��/$����ޖG���[�NNN�0����ٿ��������P5�$_G{
��?��)����M��ܔn�����ź�Ug�Ż��Cj2�m �=����뛰�c� ;;������%c+��� ����[�l#��c��l]���48��RC!�A'���W��l4��4xM��O��b)q���-�$_��?�UC%'��cu�vXk�C�Yf-8z�$�B{Y�����fӍ�.8��A�E������wC�HН�^s���#�E��e@@�� I��=b���Λ`&X$����`v��ZUѺ�N�H/_���b�iC��"�'���0iA�`�|;��@`"L��ҕ�3������٪�'��:L#��g����;(�pd�ư��n Q6��0[�b�����$c�\�M�-,j@?}}��S{j#G���^�����B�0��5 J��RVEi���g�
��&D/w4�*,��^΅w�G��~�sa)��\ ��^����%����i��w"Y�ɿ�o�m�q�
�"J���3�54��0X�V,"%��X��N���"�i�^!��c���������(�G�j��⡿&Bǹ�����rIy+b��
��z�w'�^H)X.������[�^�C�y���S��#��*Ղ�n�c;�Tʇ�O�ODy_^�.�E�vX�ʛA]_�Ϸ��Ǜ���#o���6)����+
�a���l_�U���*��^Ř'�)���{��h��"����Տ-�[@oze�J�о( �G��BB��b颥g=��޲J�6�@t՝�˩������L�q{�.�D����
=	F�0Dߤ�r��+�F���`�l;��̓%U3IM
��<��!��iR}�l>�����N]�E�H��8�"Q�� ���o��z�KyR�*��ul��5�
筝�L���ZwOw��k5N�S��*@c|- ��lyY�y�3�G��WK�qr�C_DI�����X�u��Evv���J�g����4W��8������&wv^��K�O�Aaa=X_̕A��kG��v���P*�����P�-�z�p��Q��I��#)������Qc�4��Y_Қ����bO�7�?u1��3���3S�M�i#{ۃi�<����_UTƜM�A
�.�;��T	
�)
r��D���ằ�mǜ�&n �n@\[<wi"i5�d�(�Q6z3tT�x#M�:�s
{3���o���k0�-�m��\_�.���Ġ鴎k������+�k0s��&�}|��d_�����)�l<���Hz���yy{G�����p���t�?���Y99���F}��f��v��>�������"������藧�����X�<{Ik��cH�mu��8��Ćqe�#P��[��mC��+����'u4��	L^��j�+����Գ���-Y��6�tzf+��u�X�J�s	e�砷:j�b�M��[
��
���O��]E�];�K�M��:خ2(�cVjN���5�;a�&�*F�Ɯa�؀���`��M��=�b���Z:P�s"��><���~Kn �ӊ�ШK?$�YYn�H�x�E+E�NAbj{Ϙ���g�أo<�3�K��*�I~�2�?Dm�(�ݚy�v/���Ob�6Ы��;�g���'6�2�]7xh��\�w�)+S�W.�(���@a�j�ά�;>���Of�6��gȆQ&����n���{-"ʣ $�d9����-X4H'>��H���$�w�+)7���?�s�PUkå-t�kRS}W��dnzbm�j���_T ���z����U8>/���*y5���8��uT����T�\c�q�e<�D�T�Z3��6��J1�u��wDK��ѕjT�,�c�ZM�ģ5�2�6-C�g�����
���#��3��g�s U��n`(NϝR��JnaBCA1'�E���R�O�������٘Sn:Uc��I��k�|s����	��MÜ'��a�B��:��Jd�[_��p�t�	䎲�f⤿<Yk���T��<��D����RG@蠹얕#�+~gǵ3���vs8�_�G�Ӿ��{W�����&��r(�w�u�ƈ�:(�Zy�w/x7x�\�S^��o�q�<w4}�I�2�M�����ѫ��n��2�ح��	��[��!�w�;�)+�?�I�D��1�����?�&�E> �E������q�EZ9v�fSڌ�=}C��
�&�=��
�N+R�R��g{,�%%v_�+]^� nK�=�:\CN3������'�(1)�UXukq0����r)�3-[�"L�����B�i��ة.���$���W�6�E�������>��؆ҧ	�����3-����സW8�m��0��r�V���3߂�������=�n���{JCN�d���)	���ƌ<��v͖��nR������U��Q��l���=����>��y�D�g�/y�����pA���t���*-���<_�c��>�ɐ�(�p���eR�G�y�Q��.��^ٽaU]\���RG���UO:z�d���I��#2���!�

��.耐��u^7�:U�h�X��G����ՕgN��>;)�l�-F��dw��Y��m���m�vd~�DDZ��%5�j5'���hP���wX�&dgg�JJ���V]�uk���06�-]��{��l^FU��?0)t<�ڂ�F�^�
�D�ýEI��U���V�|7O�e��<����q,H��owI3���+��sL�P7X����~�N�o�S��L��+�+}0U11��ulf�xn�����~��lF��D��{W ��yW�t�U)��e�u��:y���&��2p��or	T+s`Z��+��7��|l ����Is�f90�y�:\^��.�}������̍��ȜC����FP�/�G����O�J���	�h?��%&�����}2���N�;��JF�nť��7y��ߐ�,��kj�G>"�w�?eu�^SDKF�*^7+rc�]�]`���mO�����,��YTS�.�H���l\���>�9�{��o�k�hx�q�t�w�� �+�P�8%��gj�����$*a� Z\�T��d���=OЈfe��{	��$4�DÃ!M>�2E�d����Ql��O����9��������;9~�-.rg���g+
�Yk���f�!o����B���w����p�^t�}@�l0�����:��e?1�:h0~�I������23�@�� !���ԧ�����1�xg��+�d���١%_���:Z뷸8��[>��0D�-<�Sv�{��)k�f�.+f��X��9K�j�������wl.����)�^;��7�sy���荎�	��?mi��<�u�UVY�\Dod�N�LFTb-b�I���@"�+����7_�䣃v.�H�*D��V3n�8����9p����S�]/k�S�l��E��5�%~�/e,$�������DԿZo�i�z'�g3FG�c���Fv�o9��}��X<�y�q9&2ڤ���nk�@�dmHH�v���G&��T����+@�R�sr㒜/W��t�g���m��H�۩�x'����D�\^���o
����#�Z-Ί�u�f�b�Jx񫭽��m��}����
������P8�y�v��?��I6 �Y�wp,���Iz����8�3x21�M�,^��DS~�oo��筫�p�Ú��sI3��������ZWf��X��5lpv�L3����WT`���ͥ� "���p5�õ3��� �R�\�B�y�=PJ^^�*����}�KǗ]$K�j?��B�@a�c�8�;�����6�}`����0�en�bSãe(�o`�0 b-��o4�[�����a�1QxMU}_c.��p�,�9�����C�v����!�A��֬�i\�N/PĲ��t]: ��z(�W%��Q�����|!��wPCڂI���Rr�l����g>��9Je��N�'�4���7:7w�������uR��@��Jע�~N��I����E���G�J3�!fͼ�8���z����1�j�U�p0�ת{��ZIR�Ձ̌�.�K/؅�'G8�K�#J�^���������a	R:LB+'Q{µ|� ��$�В5:2~_QSS����IC���5B~ѫ�r���#������U�_̔W)?()�FL�.@�J=
��bG��k��g��K����<��mn��9Js��DE���	յ<+{����`���Z:kp/(���Ӌ�iF?��|��>�� ��¡FK��):��T{�4qvb��@�J��Ad>O�ձV��:�����A="fG����A
��w3~l��
e�Чq6Q]��|������3�>��P��������<����}�M�Рx�}�?Us��-�&8$�0�����D����hS�J;:��l����~�F�$�0�a��bf�$�}���pRt������w�0}Ҷ����物�1 �c�����~�u�ѳ�E��bd����yu+�><M7�42�P�+~v?nww*�D7�y<0������Nta$���1�����T�з���:����C�FJ�,�6�
mx�����(�*�/E ���6� �j��\�b�V��m�� �	4���S(%F$���*	5�Qތ���Z�m������S�����yG��_	w�&^�	��&�Y`�>��U��o����x[�x'�}���p� �a�r���n?]Ֆ�fS�uZ 0U/�L/q0�M�x��8Gq(�=�P`�,�ώ��]3\�I�ʴ�e���j����u���~��M���c�l�L9�vك�O�[F��Q:X�_�	��%'��x'�6�}��w��O��@p-�V���t��k�O��2|+?RD� ��TvK���߰vUJm-�o���� b��t�=��Δ�_|Ȝ~x7��y�x[F����I�"�'l�5��/�N����6=�]���غ؁1�v���y��zDT�M���z���4/���%�����@���F�oӧt����j)�䟠���S�w�sJ����w���'��V`�	*��}AO��ƣ�/j��R���P?1��,�.^R0��۔]T�"��HM���K9���n'��阧�R���X���1��#�kC�8O��l���.T�P��]�v|�kna���i?�	��舆1j؞�rp���a&���c	��#sT��F�
r��̼�7a��H��s�@_@��A���t��7c
T���m����n�XB3)[��d{��cZg9(�����up6�
;$�fg%<?oT�Yϑ`��
��O����)����d�K�E�o��v�Y~�������d�+�{�>_�*��$\������9���w��y	$l��T��z���:h�<�t���I�y���v@$��'�jQ��~�_�yQ�B>�M��������=G�_�K��83�V���%V����kr^a���.�������|ȭf �[����O�3�T��{�����.�#_)������}5���*��KI���c�����=�|��x���z�'c��:$;{>���Q��c����,;~�iIII%B�6PJZ��,���|��t�j�:�ʀ��K��p��gO���F)�>�6�����+�.��/-3M?ZwP ���_l`R�����֌2n�^ѓكo_�%$��H=�<jvUl��P�6}$@��?~�*�ޗn��/fDus��c����S^n��a6h �{px����M�`��,�������Y�-��3���ŉ��/X�ô^\`8���$]�5�GU�Y�� �4�X��·�y���]!���\� �ag��o�TcZtf�G���ɼ�FI?|�Ap�&�Q�2���A��LB��J�������W
�E<���:*".�c>5)1��d?�S'�Y�m����;�ay�(2��v��`���n9�xqiwH9J�k+��v;�am�(Z�t{E�կ9omݺ�]��Ivsd�ݯx�xow�y("�nG��KJB�S��F���y��\ns+�ØfU*���Wmmm=�>�M��}���[��oDuik�I��Kk'@q0	��I8y�t����jg	��qC�C�aai�!�u;�>Qlo�r�����|�?�1�B��<�xi)aKW7��XZ9��\Z��5U��ĉBE�D 0/�����\�*��@ %��������(s�<��[�4�A��IJe���o��lv[ *�!�����/�FΑP� �9���|���Nj��/~c�b�޾o]\/��'n��%����yף��!h�$4q�y@<����TR�_��f%�B���+P�2��44�a�h�Jv���s鼠wȾ��@E�q�%*�
��e+�ZAxؽ�L�y�CuA�*�)�}��#B����|Wu��	ªj2�Xw�<���Tو���2k���i���߭d���T���zp� �5_]�}�g©y���<�x)q�ڭ>��[�WΟ/�n3��!�!�>Ri�<
!����"F��yUnv���CR�n3�p�q����qP��c���fEV��RQ�Ō���9�D�� 
ō�P�ϠhђgS���a�佐�9���׼�x/k�[�x�@���X.�S,xj�
���xB��|fff[W���	�zg�����J8r�	k�o�V���Dy��3p�~h����y�O��l�"�X��8��#ǚ�PG�Pdjj���Ej��ϓ�U)u����μ��Q���(���j��W�?��	��VN/X�+�+��A����ذ���*X1�g�g�2�ӈi��E�Jxn9<��Ʉ�sy�@(\��^�W*����H��j��W�����g<~^�����"�aW-�ҨHw���*����H����.�N�����:\$�'F��O6�-��B� �����L�r�����Q
�w�t��wS�W3���$(*����>�*���y��R���9�J�'�TQ �`�ɗ��FF5�[�����O0y�z�F��A�t�DĖ��/�����w{-ܐ�Y{##�b +ߔ-+dKԋ� 6�'L��zXv����w�-SEM��r��~���k�&�b	������(��Ɣ�!�/p��	Zhb��$Vo>�̐�ˤ�*O���׮Jm�˖�۴���ta&rl���')h��u��L��ɻ~����ɽId��M��&��W�ڵo�X��b�zt��C���9�x���"ǐcuL] JT��a-W�s.��,9y�c�����O�eO�W�p�����Ap���Rү?�؍A�͖��Pn;#!툀D��#F!؟�\�$8���+n8�勯�J�)�N(�]�v_����6/�ߐ�{��>>�E[ݮ0D�,T�r���++y��}�~�i�7����j��.Cd�fK���=d]$����|����TO[\+\e~!���Q��v�E�MJ�>�#��&��g�MU���x�0W��5�P��FJPڌ ��H�|HC�{Α �@�^fm�?��hG�}6]��(P�+V6�90�҈*.�i!V�!-:�暾s�i�۾�Ģ>����x��u?7>��:�@	߆OpcB)��{�n��vA�;��f��*ټ��_�(X������!ZZ�͌�h]��5����DJe���ǆק��RW��<L�Q$ZbKVf�,P��v�z��ݤTy�Û��0t������g��O��=[����Dq��+cq�N��`~��Osn.B T��ϰ��_���2Ǌ���^����ȡ�#��8@kŢ��	ŷ�~��o9)�0\(޵����} 29�}/-ō�}�6�#5t����ǹuv� B�R*w����@gSӤ���l�E�X��2wڵh��¹u~_\�W���莂[*�Qy�vm}�q�d�0����&.44�2ؒ�7�r�����a+y�SS
.�ɼ7��A���ѓ�_��j�Oh�L��5��^O����JALT&U����1f��p<�O�|Y�����R�,���Mc�]{���3���U��T����A���,���4��e(Q]�V]x���0��]�\m+S�+|ڠy�Bkҏ�^��^� _�p����bA?�M�7
ơ�.�����
 �1��B�U�D��66&�6�I��qe,F��,����(���Y
D��ظd�dc��D�����]o�U����P'��(̀��s��ڑ˱;��.D�ܴ�$�§���n=���h0��s����#��O<>n��j-R��ۦ�X�#^��s�l��_%5��ş��95'���";�GjpLJ���ɿjW����p��y�&�A+�؀�����kW1[��A,z��v 1��=�TqS�!��I[kf��(��{_���(�%�mѩ��<��1��C!k���߁)p[�()��'Dΰ��/��=��j��~� ��>�\�o+;̬=� "L�w��RQᴩ���|��V��s��>�W����������h��p���C@�^�0[�.����c-�E�+V�uT�;�`r_K��OK�kNe����̡�£}$��=Qf֙�6Or8���r�,;/���Z�h�K?�������A���s
��������ׄ��߻��#�P,��l�ΰ0�P~%�#�4un{�a�>�c���2c0�6�#��ї.��=���ɑ��xV(sA��TË�O�b�Ϫ��h^�?��͂kv���g �+*F��L<h��G����u�^��	777��`���e��_��<����tXR��"I%|�>����l�w}K`#_�U����y���N/b���Dr�I}���*��|�'%�OJ�;0��2�|"���bO�+���J	9��U�J�OR�.��j� �`l���v�CB��mR����_Ǖ��q��%
'��T�"Y�nUQ�d^O��-P�#7V.�bW�Vk\���D�J+�;����u�7!l���Y	�cՂ�B�X\r\�K�^��'IA%ѯU�#��w����%��_��-I�h�_&���ɓ��p-k��D���e���C���l����3Z+�:���㱐[tN[�&���i㌣Mjƭ��Kd��DG<o���������\w%:�v
才�k}Y�a ��xU��QV,��HF�zC$�i��\6j�;�����8
]�c�?ڃ�i�:!���OM���\��4�L)L��O�T1 ��g����)PYq&�s��ͦ��@�y��h������+�����{��&��6q�i��ۋ�I|���������t{���$�V��Z�6���Of�^PhlqE
kM��0[�E8>(ܖ�z�6�"��$.DU]������B��a����gjhr�yI[+,GB�{��6E��NL13p�� ���Z�����|�Mr�q���E�͓B�K;�B�'��q[�����r�����(�VoN��"}
��~~�M+d����O����Df�􉂱�Z����`S'��K�'�f�=[!�%���/�!h;Q���2"<����m?⼣@�Й���WS�Ren�Ω�vrgL��$'�0�#�Z�3bmT����Hwj��kl�үG��	_6x�.w7U{G-Q�(� �b13�&y`N��1���!P��G�J�>_=�������˾ⓗdx����r�G����bani��;_����&e�
�^�5c�cN�
$�yǏ�G���,?���)p�;���?�[$�
��}SR2�����U9��+LTjU�ZW����m�+j��@��y�I6V�ܙ��1�D�=z~~~�G��ju����YH!�[d3��V�V�A��}����˰�1��J�w�_ܻwܿ��߁t�f\����t9��X�OO��}�oÈ�"<�M�K�xuI�Mc�d��3��޿Zbm����_̫1���� sӕ�~|��^��|�X��C�x���JTi����3*y)�w�yg��������h"bg�X�����W�V�L�nֺ4h���\�3E���^g �9�jg�!W/.��	B>�ȿu�׉�>�A�-�mKe�>��g�6`��LN�3�`�+n��qʷ��W�V��0�q�*t���z��,��I؏��V{�,"?�\i����W��H����T&X�Y�]޿�.�;5�q4,L=��\��R���n��uo��h�;��A��3[Vጩ@�hfY�v��(v�8�.�g��5���?yv��=s��0~.G�XõuMѱGl09"V��
��4��+uǌ@�>�
4Uut��D�_�;o�?�Npio��s\OOq�oa鄪WA�J#i�俚�v��ҽ>�۪��$;qO\?*� �e-)�g��Y_�3o��m�un'�4.x$�ɟH�R6�=[�<���H��<}��{M_v�@!�ϛ�[|(�#����g�AKA���Ǉ��5��g�$��D��4���/w8�딸�El��,�+���y��S�$:�y�t�nu� �'���F���"�c�tș��	���3�ۿٴ�B��og��_�豮�h�����*#�[ӯ�P����2��|��=ެ��������ϗ�z=���o��l�1�-�.&:�H�Ȩ�|���J��Z�j�/����/�./G��K�ETQ��vO
�G�϶�B���]�l��N��o�Syi{˲�J���;��sz4��9���cټ�MZl?h��|��)����1D� ������(��Ir�CII�}l.��&�7���X*}�WK4|�`b��P[�&��|Fj�ɖ�&��o��b�z^Vx���N�.�k�Ya�.���qӎi���G�������Xw/�z�>%T�\��Y�W�=�[��6�Z��0K�3���M���x����[/��F{�i-�� ����g}�
d@����X��(,�"��I�d��Gr}����`|X��_� X��/����)���zu���X���|���!r���(ψ��C�S�! 4�[�)l�T6A���@k���8K�iCgDr_�Dw�<���� ��WEo��"�E���b�$��J��e��w.[N�U1�T��xr�{�b��u�Bb%`K��j�9���i5��¿ #�@Yv�67?5�VT��	`��A��K@Ka2���H�9ٙ}c����AO�-^ty��y1���j����Gڴ�?1�Yا�
��+hf���b��n�T��h�|/C��z�Ɨ�ଃ���R��=��{f�{9�D�����!��`A]Թ*Q6�#i4]ٺc:7E�=w(e��3��}��B��$7�´zb�c�0���f3P['q�u�(��l�:�G�e�����p�G>Q��J����E_˵�ļ:x�Gz׾�Ϋ�2���p4�֌���`�џg��y��p��QKg4��7wu.�OpǺnF�G����(���}��k4Re��uka��{ޕ�:<;uM��e� Ck��A�W�"@�w&�H �U��%��$�{cg�)Ik\�ׯV>���'ʪH����oM��Q��k�>��{\�W�v~�;�:kLs��b�/�T�C`ؚ�Pa
�����H�n����hL��y��k��S}��97m��k�ϊ�� yl�e��l�I������$�+����_6���˞��},�n���#��r�u��>��g�b:�eq��Fc4�h� 5#4*t�ll��([?�[f�)aCq:����[����ـ���m�9]�Pm���ٿ���O��bW�|_��s���|��Hy�\�ܶGs��-���TՀ������}�����%��9O���K��K���(��|��$X@ƙe���a�"w;�"o��o��Ke������n8��Vf��"�O>vC�j*0��h�����ᄭ|60�O%L��Yn�_m�c��"W������{9nz9�R�H���YL��<V��M�B:��x�//��z�;o�M��6��h��]��M�N~���g��u0y����5`7��bg�����r��ѧo���f�hj�&�:3p�����&����"��)�X�H �"ɦ;�3/�Gb(O�%Ѧ��a���)[���ȳ��!�&�X�M��%PY��g��w�>��.�QSz�㧢Ec�j��	�H2.�O�S�g��Hq�*#�A��(��'M�Tx��L<�Zz�	dbP'���?}���Ŋ�SLRw.0��1=z��ʡ7	ﺻ����2���wD����}��X�f����xx}͋���"��»KA�y=I5e����z��g3f/�i���Qg�M�=����.�0)��a�߶�A�6ZzR(���c1-�uA��|��Ϗ��ú�?j�x��%j�x������307'��f�+�H��枿62Ҥ��>�V[�#''g�9��p�q�L��5F4��Nh�&��~�.߫zI�	���G˸��bW�*��$��{�_:����g�5#{�*Q�#��z�Ol���M�q� Wx�W���Ee �!�����Z�Y5̆��ﶸ�V�G߂���
��n�z��}���	[�J~�(o˵���7gpw����-[��ڎQVLX*�k/6`-���
M]}ǭ6���:D&D�0�p��H���������ނ�g���A�+\�����L8N�\�!nZ:��@#�R�C�����/��Kc��(�Mhk�\�����W��k�~id*�M�-�|��}1����{�R�k�����KUv^�QN�D�cA5���ҟ =-*b�iO:r���=6#٤\K��E������'�A��-���X�����է#\�����ܱ�rIءD�d|`9�p�JuRx�}\����6�ɗ+�ۙ��{´ztD�zȈ��B�UzK����칈ݦev��h�v�#:[�;���E*yoL��ȉ��U
<oc��2N��1m��q�@(>�����f�I0]�<;��/��1���@�S�"�?�߈g&�႖�9#�1���G�d�:�c�M��'�����K)Qbb'�����8�gv$6&A��E`�U&)�z�Sc�3��������ĥp�T���R@��װؘxO��rm1��!>�|y�������u���{��_
c& ׭�K�|Z;N�x8�)������s-Q[���;<��5W����b���-�Ğ�viK����nsrrzU?c���8��](���k��m_�5"VJ뜱D�oqsju/������w��?��w�����}�ٙ&u�&X^ɰ����X��8�+�e��_6ƚ�2Eb���Y�g�vlf��$��#�m��B��T�򆾧����J7D�W$�#p ��"�3�|�b�]!��-Z�c�fQ����c;�y[/גV[��ٕ6����������o�:c�"/�-A�Y�t;2��C<XӁo&p_(�������⾁��SQ��T����rHR��[s��uu4����!6X^-
sL�|�wmWgq����ay��q��F��u���a�m>>�Hl���W�?ջ���w�ΌC�N�\���*վ��f�P�0pa��s�r�ح� ����)s�\Z;iy��z���O��wmZQ�?WNYcm��m�J81a��煺�f)��V����� �7�wT�hy>����_��b��$	J�����K�_p^�@�ZD���mպ�]��4r�R53s ����/�������h�|Ѣ&+>�:3��I����$���Q�M�l���<��[%@��f`�K����C��9r���ʨ�x���R3	aP-�^.;����_���=G`1�͜�O�U�j+�����PmvK�4`-�	�ݑ���ڕ�������_$�,��:��ц1E�_y'ݞ�ˡR%ʖyx��G�q��K��s��H�h��4v> �V<�/�{qQ�z��{~�����10�'|wWv�@�j���Z�����k���m}�o��=D�&M?���Ryat����;������U1��l��Z��鬧u[�]�̫���`Mԓd�<�1)(����y�<пg"����OA�d�		 O�|�Et0?�{.�'���?��d��W�l<<LQ��J�=�+i?;+��8��i����g�Z�a�]�Z:fh���Y\[����]�H8����,�[���8�t��I+�߿.�qO���>�̳�]V���=�P(|>�#���y;��՛�4��ݏl�y��K0I�FFf�P�9��Q\�E�ɍz����:B���Z���$��w��K����=a+g�	��`ǆ�T�Hę4��7Sd�1>�I�Іu�+�V=ދ�p	�Ķ�!W�[���w�tI�7�A�ZGJ�4���%�[%��sp��H�����w[̜e�t%wĿ����`(����.�]�u��t+>_qb��J�����H|�T���l��V�9�nA�ʽ���ؖ1������N�?J�(���F�Mt�l4UK�(޸&�Q|k�|h�rX`��=�Ժo��)y�Gj�-�t�y`���(����M�n��3��S�y��՞���%
����U�9b͎�"I�5y��5\|�$����DJ#��]�?D(
w4�("#q�G?�*p+w,��-�oK���W���K�<���&�zlQ��g�H����V��ߊ��f�c��2�g8�w�ӎ�=3��<�2ؾb�b�&�jp�&N�F%d0�[�e�=ߜ�4���a�����Ӟh>o�ڪ+�t3�4\H!��z;_�v�j���|�C DK�j�ms^��c�""�U�O'��,~/�7}��$=����-�ں��1-ew��w[בq�����K��J�+���(�!ytTg�<�����ٵ����pp�H��	��`��׹�X|�����Q_k�����7u�x��g��4���}��G_���(�`��$.�=M�}lus�kniiN����n��N\m�_��60�Ä�tN7xabc���hy��#�X\���WX)��0�sP$��Yh��*�U���S�zOl���.:��d	'�����g��"ma��/lk�h�PI�P�tJ�g�NO.���EPM�ߓ ���v�t���c��	�{�>G&���o)d��p1�I�o^�!��Ş�}� P������03<Yn╛��u��l�������Ѣ�f�X��*j���(j�U�*j��j�V՞U�Mլj��?���{���{ν�����y���uM�v@�޿���X�Fb7�8�rvϚ"}���x_�E�f%l�gJ��~X�<�sU�!Z6rN�R|��M���~1����~��2u:n��M���y�fbYRV�I��Mc(��oB��w��J���"�M��Ƙ�_�ۺ��}naf��Ԃ��HQ��cKt9><d/��oD"�v:�p�ՆVȯb_��
�N�TUs�	�P��%$����꠻��)�V�Qlͫ@�tg[�>�[�U���
�f|+��<��Z���
N�O$�,$ɰ��!E4��@�>��{��XhNNk��G{]�N5���k)J����l��Y�׷���>^���|����[E���R�猝�������=�����P2��9\�4�z��\�z@)� �}R&.,l޻\(��Y�����5�����v�߉���;j�?Y��1����'TCM8��#M79<z�h�V2��$,W��/'mopS�}�. �ߘW�i;�=�g��||r0[���*TO��F�k�BY�U!Ѵ��O;+βT���a�|q�U�B��S��x�R��uP{�E6��o���H���<A�[+�thzNoW�.��O��)��[+}��y�ԯЀk,06l�h!S��+�Y��&G��wl����ۧ�Z�*�L�+|}v��Jt(�W0+�G6;e��d�t:��*����������P[�/Pc�f\ǈRXC�3�U��yQ'Wh=�?�<�PT���MF����*�io>�cP�p�8��_g)�r}/,�h陡�&��̙e<Eu�tt�pV��J��HW����Q��a����&ƙO�7F�Ytp�AN��E�9h�B�D�}��	�wg���H괌v黻+���'��]��6��17%��S#	���ۤQ�+�ek3��>�~�dq��asRT6?5Yh _s\aJ�n�{�N� �֜Tn��`����i*dO��bj�ǉ�9��7�]���+N��������ص�����us�I"^�H�bT��T?S�K6��˱�����8K�oN�A4��c�M����q`�W��o?�ؑ�9���G���J�n��͎C�ˇ�;��RM�HW��|�������)0ɼ㡁��g����!Pj\S��?�˟�s�������d$xn?eƲfY3�P5Ҩ�|{K��B��1;�X��ut�'�nb�:A��9-���������]m������d�J��WE;#>U�O]��\�g�������DO8�	<\�>�3NHQxҭ�8�fH��o���9����(V�]�^�%'���^}MR��qA]�,����A]=?�Lh0��I��h��Z<Z�o�F�5E��FZؙ��L��	S�>�����*�-�~�:�W�0o6�|-o%���*�����Ә�����_�[��oDl��zm�t�p��>y��>� �IN�y���:�=�\N�?C��)3Jy�-���&����������Ht��X�)�Rx1a��_���dY�q���+����q;�)�U�w\}
G�?[^`e�n���o�.�=��fC����0bO�S��݅1�A�4�#���d�����&1�g�%��G��o��e'@#��4�H��g=<QCfn���ʳ����^[_����s}(u�`�	�/�^59z[�^�w&�|R�;��N��\Xi�F��u�~��!6�%���sd�L�V��)+�̃H������
��n�=M/��<ߩ}SV��b���O� -ډ�uKfeO��8��8��5\��s�+��5��W�0��0 ԌtTFR���W��4��Ŗqv��k�&��p�K��f`�7Ó�7�(��5R}F,:�F�V76�sЙNI(��N.jn�ᣢqQ��1TFC��ߘ� �D�Q8MO��=��q�_uBu0�$�4�AN�e����ʔ:���:+!ԅA�31ˍ'6��U7W59��W��)��j���2y�;�L2�!��?�"��*}�����}��YK��6�u7򶰅y�&a��̳߻?3N�l\��HXC��ya������R�&{��X�aɁ��.��3����#Q�y9N�������k.-��	�kzPg�IݥY�����	�'�����5(>�'�+�l�o��Y�Uԟm9p�!M�_8��C��Z�Y�v=?KR�k�D[j`q��/b8��E����{m�@2X����xзf�����Ad��u�g� Tf���}�jrɮ*MjS^�
#wZ�W�wȮ�C7�ME>���H�'=�r��A޽��s��D�-��P�~Y��Q�
��BqO�ba�N�@�-ݢfo�TZ6�ί$zƧX^�b�nL/�?��&P��`�=OG��;횃�M� ���}�{V�}a7b`&���yq�h{s��5�a�Ԗ�)9y��%l� ����.3�m�M��݋�������'j��\��-@�ǉ�7��H&g^��\��BVw?P��3(����?��h>��-�ue��ķ8Y3��C�ge��f�b��� %�)�ĭ�n�k9��fk J�:�v1�n�t�c��xX���?q�u"<΅g��gP�JH�IduxG>(�QW`zu��L�����@��3Π��	v�P�/���js��/��ų�nUx\otv����o����Qډ��b?䐐�V`��X�h`*ؼ�'���J��s�3��#�\O�na@��14P��تL�0@S=���l%��j!n������ P����B���9���S�ׂfI���z$\���M>��)���/hcY3��И�c�&Z]C�����u������M�s�����b��d�E�a�h�G>��vҚ9��7ݿJ6{���+,NY�򵕪�I ��wq���D�r�r��u��k6���v��v�:imH�B c$�}J�3������w8����4o�F���b3!0�\sBPğS[�P����V�=�N��MÀ����[�}�N[���|&|�9�����JUYݽ
ɩ�LX�6�9�����6�Ԯ+�i��;�idI���L�l3YJ.�����R���zP��d��Xk��Eƽck��������1�qN@�8��w�R��#�9����B�V�����W��|���:��f`M���ʀ�|���0����Ͷ���h\�x�� �6���܅#Y����ϗ���SZ���S�,����	�0yܸ������k(��6�6n���&���i��|�>Z�׳�~�f�+���Om�p�o���:S��F�t���?�vXe�(a�Z����N�w	#c��A��2v�|=��N .V�$[;?�1�LSF�f��A�c��d�v���h����'���$��w.%��[���W��\N�0\b�(ڽ�:�����nu�#I@8C�a�8k�ʉZ�]Ȳ1Ϥ�� YB��Dk}��Y�#eJV��. ��sP�!�V����X�%�	�v�eԒ�����+s��b@tȮ�p�j���K����J���9�e��oGM�'<Iq�<^�6qo�jI�Ã�	�+��5e�� 0�*��ޑc�
�[0���5���Gw);0VU�߭��!r�E�i�@ X}�Bg�g��LxX�y��a���K�G���Sǐ�����b���Zf���l�q����r���b�᧱Ͱ[���Wy��"������t�������y�u��C����/�?�P�2[��_k_�2<*#�wv���7��p\��ww�.�C��dI�G����'�>�/�^8�4FkM�`�3��;Ӏ���=��-�e�ɘ��6�QKl��*�̒[���ѡ��?ﳵ��d�W)�D�����$!����=[�&�0fȧ�{��+Lz:�F>�.*���bq���I�i8��u�����,;��ɉ�G��������N�n��-Լ �,�*��^�~�]�s��%Hì.B�(�PIMW>�gQ4:��*�X�K���
��/����/�q���`��T�d"�Բ%�A�K�>�hN��M&� ��ِ���͉�gCd8!�d-!!!�CL��J�Z��ֈ��0qY2��t������[�E�O���������'�Z���Ds)nx��H�	1`'���N��=8�+�,��*�����REH>��Y����Z|�#�\�� �ٽ���K�K*��xcSW���{���0	�U
<�\����~�+���(��Ù�B]�籡������Td�j�;�\��K��k?\�_'S�z��zaf�_O:�-1ZW��l��$��A���@T��1�e��}���m��.䮙���@�n�_
�%ף$?�����L
UU�����Mt���\���o����9�\ on�����/�1��aq�-2����Bi�qq��;��?"���F�M	�$�[�rI��;Qļ7�3�]�1\ZL��V���˾����w[Pi����թ�[P�8�h��Ad��
V��p���E�R�~��/�z��1���r�m�j.}N�1�|�{���3
�è�"��7������zͼ�Ԛ����O1J8~7_��wwY�O�Y�n8S��<�>;s�?�y���ɯO{B��c��?XjO�UEˊ�)��7�$E-/��K��1�b���Q�(QL5��		l�q��H%�z]}܂��A���k׮[~�τs����	���t�υ�5v
΀%�N����gO�<��T��k�
�t?y@3%nÕ��8�|��Ł19�3��T�̶�0��Ānۗ�j��х�U�!5�{�&L�
����~�&2 Aŋ0��]�������Z6��5�'��4���7�@,B�[�0�Q��z�`�T�B�'���D<ܖ����c�T�BZ��-�� ��
Lz�*L���H?�!ωE���TX~���H;���2s),�P���nԖ�� �Ͳ[�Y�WLPa*�L?`,Ph�|T�:�bg����QxRևH~в@��~�C�x�^�!���J�l�a��!�,㴌��DJo��>�q`j� ���V�܁;�sj	�Qj�O=3dl�JT^�x����K��ڟ1����)��!��N��2,�sIUk&~�#�4e#�0�stҞr��pR��4@������YS8Ѳ~@c��rB�\��ֈ�d.��Ƒ��@���2C>��C%��C�	��G���5�y��~.����>�3wia����a�!���}26���$����Ue�w?
,By�d(L���:��S⽖�F��v���%,�uK2~��Ɲ�^'$��bV�d��0�%�I.dkV�Y�O��Kf�#0�Ac��݂���FF�^x�xT����+4p/.}�ּ�ҼУ��Y�?^V���k���'WW��KxRMb����ϳ�n��Ll��X��M�F�6i-��T\�4oa͎T��Z�"Rȩ���h�O־\�X��_;��W��������kׯ�7�-�\�n}Y�V�sX�|@��������|c~#����|�Η�ѩ���v��JͿ���%�3EfҐ�Y�Vsʭ��u��:�������w�J6�ܡ��l
���u�Rzب��Ds��[E���ɤ��f��%�vG7��W�A���e�����������_����t�SA �{��a��P�uΜ2�>
��%w����(D�=���v��|\��	"h���u�����A��̮|
X��A�Vf�z��A��������8�����B��zo�{k~��>�=H�4J�K�
j��AH*�#��������Gj��7��w�u���&$r|�xǩ�HX�K����D߷��q�ec����`W�cH	�����9�p�%	+U���yL�i���zקN	�{H�_V�������ghMHZfږ�\~!O*��[y��`b���[?�y�1C�m��`�Ⱦ$��H�,���6f�ّ3��>A��?~,��.v݄Ɩ﹢i+R�)ǚ����\-K��F~�'}�dyiAՆ�[��:�b+ �[Q�[[���Z'!ԡ�>�������w����r T�;�7+X��A	�
L�2<P�qv1}�˚���}�;ӝH�� '#�	����t�����|\)P��_��aI0�� ��G��U�*X�TX����u��Q���{E�v��*-V.�z{����M�=8�|ph4���LNGg�SқW3��J9=�͡�O`��LH���%��ou�L�e�����u��6/Q�sf[H����b���IƘ6�N��s=�q����;�|�93-�6��M9�u ~����x6i��NA��XO⼏J�9��]�(���(Y?�Y}:|�<�4=gP�v��a���E$�k0����K+ꮍa_��\���w.���=���]U^����>3�=ǋ�G���G�w���u�喑ۖ��r�hD�oB3G=��$����n8���ޭ��� %`0:�5b0�L�~��N��@oxHS$���i�����_A�� ȃ��Nx��Z��ă"�TVV�iNƏU��$�T���-m�M�����j~�d��|ŭ�{���޼no�����8����k!N5[9xXcJ��nX�-��F�����e�׽��/+c�>v�r5�F_�|Lu+H�W�k�8�L��?c����]�ia*�a��'�rh�J�@�ԛ�T�)�WO�\��8K�ph3he]��&o8WсUo�wZg=%��T�/��'�ũ�JHv	&Ő���k���\)�cݦ�g�ۀ�;���י�.�(cȲ�09��Hl͋ܵ��KS`2�^��(�y��7�E���A�T�������^ �շ����w����ٳ�{ �� A�Mс��zS{�� }_�Ug*��]=8�l���8��d�	�nz���Q5GN�χ ����j�󔉗��
 t_�+<6�r�JU�������,Ux��'����p[e3���o�����~k�R|o�����7���%e����eU�L<T��`������!+K�E�v�£U��c^�_�1�"���W,��� r��)h��[���
�d����hy���!=y���p�t�-v������s-*�z#m:��	�|Q0z��8���&ϕ�;��\�� �������GU�:J2���g�eD�OV+�vg�7KIHPWWzQ�!d�o����^d�Vk�MNf]%�#����ԕ^4��������\�2>~�J��0�6�4�9o�������d�싞J�*���W�2tm��H�P�f�[��oZ��$*(L�Kl�0 3׌S��r̟o݆����/��&łR�5�#S�����،��6L�n���wj���hZTT���]U��j��?n���,�y��K���g�S~�� �ڟf������3d�UR���ݿ�����lޅ=�T_������`�!ǯ���<�25���H��\��<X�iZ�'������r��~Xz��֟�<���6���v�MO'��;�i2���X�=���P������d���aas�:�@�er$�3C.K����q��o%L��O���.�Ur�����խ-�T���T��@oV�/#�ùm�4�������K6��
J�Gt�qƟ^�}�g?���ނP�Ó�M��G�lv�m�+1r�
ց�L��i��@�oR���gMu揈��8�eU �̉p��F�����	�x�_t4�y�T���RA����|���:�1j�qo�C�(	A�Ň$"-H�N7����W�����-�$BW�����8˰���]>��9ef��k31�~�?�N�}M>ֈ?��I^�]m]`>%��	7�ÿ���������oi���y`	�.HU���	X��dܜ�'V+U�H�$bZ��˟�;8�$<��|~�/��7kAM�]pT�uP.���o���J�����5y�i��x�i}i_ӕ, �I�}���w�n�m��܌��<�H*]��]�,m�7�K� �x�"P-�d��>���1�d�(R�+��w�P�õ�U�����e��]���*����-���93	֥}$b&``ʫU��7�y��gVe����Տ��k*U`VD�bL=2��˙�̘>̉=�d�B����*�!�:��7�Ё[�B��4��J��3r��?#�q��~�`9`��M	��s5I��3D&�͠���&Vʔ&hcOB-���l�)2i�J|��Kz��~ωPh6��F�/��F�q8_�[�N�L�� �t�_��CB�XG`�x��%���A�?��%��FKJn��YY���z������A��ib�m�ٓ�{��z���<l��q* �cry�-C��\��	wj϶{��P���+�o�� %�q����çR�.C���-�' MQoo�<=��~o�~Ⱥ�c��7J���N朶�x�W`R,��ޫ� �I���9$������d�}m`
ɔ��mT{�ddp��B�}xCC#�j0��q�:��fH7��<H�ܥ#ɟ�����x��%�~o/�FwN"�$R�ɝ�y�=g�[~)����%�|�!OS"��oIQy�`fR���l���#��b. Ŕ�����д�J���I�*��z��C�D��B�W���>.��&��$�e�U��h�+��ޣ��O�:�,�0m���t�.W����ڏ���\?�Y՞��w̕�(��e��`��*�0���r�oN68?��U�8����Թ(�Үw�AQ�u}���[�nXe6t�C�m�0�i�8���Z�Ϊ+�,�+W��V�?mȍ��� �c��I�k���v������Z�(����X�Ot�#I\7.A|��J���1���M��}q� 	��x5t����hж�0d���'�5E�fg�X�/C��`6K�C�~���DP�B.gʻsQ���[H�=\/�*�tu��!_�y^wգj���ӻHhEV�o>)aVK���,�!&�_L1�>���h�����E,B�ק�(JM�!���R�>�U�"�-�ب��M8e"당��J#w��܃0���]�Վ�� �9��ƞ�����v����g��f�a���U=X9(u�rp���d����&��~�k2����0�׊ic�$�leޛ���xO�Տd���휌O�����LLM{��d��	�1q��}O��	+M����IY<E�^dc�?�e�~̃�o����yxZ-^ �d���0"}g�%�̂I�\�va��B+��y����� 1�;�nhzZ�I(�ȺS=�N�|��1/D��5��r��~23/+�z9]�P�2�.do	�b�S��f@`��!����K�7��4��T@��.-U�����  R�Cv�	�/bD�"���[/.��<�>k�BU�mS��hn� Kc�u�o �pw�N�a_^���6!�(
		]5�4��+N��H����Z��q��������'fwB�S�撾��,�;� �#<�t*����O>l4�Uh�՞��2�-�|��M���$&+��
)`�O��f�������.Z�+�q�^��H���,:YQ˴/-pb%�©W?W.'z�_<��k��%�:372�b���׬1_{[��9����������ԋGZh	�>��Uy�͍-u��z�q��XD!6��B-)V� ��c�%Q�`�w��+q�����a�e��O[+^�-� �W�e�z8��O�C3C�4�,��1�S�f��Z�3�����`�& z�%�z[�m_Qh�SH��w��@N��a^� ��h�!Z2"�!���>��D���X��;��f����8����9�ȝa}��H�[!�t��B*�;eo��]���b@,�Û��� ��-�Fu��S�Ș��p�����Gnl���"���.�������'�nOE8�Z��"�z.�=R��e��C$��$yR�� '@2�(Ɋ86q�[R`�s��d ����z��Q��4�fL�	�z��A5jY�w3$���A����bu	w�g�ࢣo�D���4�h���&:"f>ް�*D3�`�Hw�/m"��FL�Ζ�5��ة����
w��;�ϻ�IHV��BIfy�|s��>���O�xu���Mf�K����8>.(�Ӂ7��\ ib*1�ľ�.v*�k;�u$��-	\��唯�]-G���H����� �1_GB��rʚZ���a�U���d�$V����WXVUa9ԥ������`��l"J|�_�p��q\¾����P�����>2����n��h��+Yݗ�=F��BXՁ��Am-C��(Y��$ՙ�b+��s����y����p���VAK�%��<f>rx����-}�qh��3�4O�"x�G�Uq� 5G��X#W�y�\}}Q��"�f\��_ɏ�td~R,k x]\�~)��n��!&ߜ�`�w.�1'8٢5��mU�E�z_���נ��P��#��	�p+�2�7�[b��/�p;Y��hs�Ĵ[���L��kA�7���+ �Uc���_S�vMo��ܪV��Q_����PR�O�Y��f��~z�5G����	9z��2l�oӇqTU�@2�P��%	��}!��,Ӡ8
��)�����3��o��i��xԴ� ��9-�*���/�X�EL62��x*�d�=��/���=��VIŸAԢ_�$GG��Z49��#�۔<�v�5�FZ$��;sx;��p��;�i�Sϣ�t�_���c�7�;΢�,�!4�3��u��
9,��i����c�&���IȲ�W��1l��G���e Y��k�iJ�-Q��iG9x�Ө���^U�O�xI��J���F8C��>�Sm�驲ٳ�����Q���)b���XU�j~�x��z�����c-�Y4]:
��5�!|��*k��^�S��ڝ��='c��q�u�\��SM�+	����\
�$J�;�eP4�|F�P7��-�~e��oX��oA_g�F5NL�ڕ͘X,��{N����OU ty_��!��ю���>b6Em:���7����"J�ӎo>S7;�o!5������}��������]w#�?���d�<�`doW"����׭����Vw�v&��w8���/����W)�q,�99�s�AW'�s?uuqy��)N�*j��n���X����r�;\�^�y�=���:��1O�tɓ�u����8�WlR������d��P@��(6��Jx�0_��)���I��|i {��¤_%kě�� R�T�Tx��0�!��8�~��������8	�l?�D\�D�N�j}���H����o��𰑟�]$���k/�H�4��N��nF�R�U�࿹ �/����(q����L��HY���NEV"�x���G�>($�W\'�C6�yH��3;�lXڻ�\Ʃi���TL�/�ޚ�'� *Hl�'1�1X+�w5uD�)�/�nMŚ�Z
����dY��RQ�iu*4K�8�6C�k\�ɯ�O��T����Z�|s�j��N�kL���Q�˶A@W��5�*n#��R��(bܞ]����	��
��Yx-��ج��B�I1�%v��䝟�.*�H�j�k�27@�XOcW��;ot�,x�n�G��BhL�G�	3C���|��8{��vmX�,��+���ӽ�!��N����f!�/�3z�����1�3%���w�b�51J"L�s�b'��{�80)��5�TQ}������r��rA��i=0��ζ�A����#0Hَ�@2t}���~������K=4��W�*�(���dJ5N�]���2 �����!֞O�@ٯd:�9C�>�0�ߺ�n{ש�̝2��Ձ����M�U���f�
�N�t�t����(��X0�)�;o^,���/����)�����3��N~�5:###`�p.��x(��#�"��6�m�j�f�Ez��w.h��l�]�:���
Bs&��ݔ�<�7��PP�Ǝ������dy�"u,+�.����T2��-�xv�@�g�%wh��Z͐���P��	�[��#;f��-���Y��2a��I�uV+q=�O��A�f��++�?T5��yMV\��$Z���u�:#�߾����Qw
�:�z$�a�����J1J����]I�/ *��KQ7�FW���5Qh����ٷ]�a��Q��+JzZ_�:'/����+�4[���m�B�UH�\OY-�_�l��Q�/��.�R�e!���_���ɱ4VF�)��^���P�@�W�qI��Q�[-Qc����6#����3�Y��xۈ�t����&2�����}��K��^Ā��n\���x��~b���yG$rK�q�pq] 6#E͂-}� ��[���3j�.6�z�;@F�R'��b��{����4Ɲ�@�zRj�L��@V`�F�!$
�_园��q�H('��c�_��Y��� 0�e|�]G������,F��&n�(�[7�p�[wo���?$����Ǘ�M�;��SdS)��� �S�L���L���Z6U�*[ �������1�O�wx��)����*�όx1�	x�`��U^����Y�R=�6��O^n�eqb�=��\u{#'�#����Y�b�u���K�*F��������B�fu�׷�^��ƕ��=W�O�~�1d���}a�DFK�p׆�ҏ|3׮�)�k
���:�ϊ���P�|l͙=�޶q/���K&o���Á�n;0�C.x8<�{�Gi	�s�AY���oM4�G��T�z��zN��0��rc#)*:��≚
;Tq��]?	�������rDX7�Z�j�ꇟ1�v*���Μ�0	�
��d�U���y��WJݘT*q�ْ��ߨzQpc5_b;��[����Ub9"٩k���l��Wv_�����ϩ���ڛϜ���D�T�t�����qɴc*%�^W2�m=O �WQ�v��	��+K{F���m�w�u��Oh9�r�J���F��fq�X� ��$�ɭP}K�6�9�#1e?G��ތѣ����슧�#��n��Ӯߵ��G��T3��Y�#�.�
�r�M1�ێ�����v_�')�0�Ϲ\��� U�	�ѹ��Q����D���QF�@X���3&��`�<#�p]J�̽����(��>Z��ɺb"tA��`��l��U�T7����U)�hH����°X\�h���!���?Zf�1�
���?Y��EMY�_y�����=M�$hU�5���$Q4���A�?SeRs5KS�*@I�S>0x����71a3�Ϸ�(�9��[?"�n�C�������T��h�Hy^��Y1y�T?i Վaw~/���2��6�vRh&�Wm6$��W0MC�J�������ճ}��8ʝT�(F���fmR��4,�O���}*�b�es�ܣS���|{���SM �~��r�+�� �q˔�kVjX�Z"6��7������%u���U������M��>��G�c���dHJA;�Wv�8�=]�VC4Ww�w:�^��}A}�\�;<������2%L�V���1
:*#^���t���G����-��к��	�O��P7&a_��[)�%�y
l�"J�>T~�ڄ�:�CP$��0���Ak��Ǳ"?��X��9��P����4��0)�apf��80����I�H���P$ŤO��-�~p߭�rB�I&�kR7o���k���;jy-\���RF��=-!\X�/���&� �����{���Q�^�J���jb	�8?������A �����qǈZ�^�w����8K�w��K�mTII����u>K2%ۻ�]s�;ƀ(t"<tk��������e�e���B��S����/4�m���r����������m[] 7������b�����lB���z]�@U���Y}E�+,���G�npc�#�Лj�����޲�Fd�%BetPyJ-C��QcJO/h
G|nUdƕ3E�H���P[D"X���?� H����C!�Z��Z�[�/����[�]
x�[�&R,24�ڗ���L��i�ͷ%b��9����L5��aH�5�Ʈ�T6�C�vlq'�i�����s2����*-�����>���Q�҆�٨�@ȡ"6��!��~0�z��y,0#r��F-�Ց�Sî6���r3m�f��ɧ�%/�ME㡽Q���9X�#M/;ZX���ۥ� �ؑݎL[�T�D��'r�qg�Ί��5�K�Go֣�*M�����K��܁7�0��K��V�K&Nv�O���n�_w4�Ե�g���r�L�W�Y�pq���E�Q����2cm�k@�������=BM�i�;�Z��n�w	�5�y#��c5�d����U���r�����A)��zO��7q�i��,&h�O�b0w
��3q����I�ؙ3�:r�2lRq�tP������+�7qCsH�񀩳���O]Χ������$�����^''�R,�:��Ņ�P�`4c.|�$L@�����ң}\�N�	4�蒾�2��_C��J�_H0W�N���q�LI�] ���B��C�qX�����{�/K/�Y�<xN��������屖��G/��?�'����7T,	!8}_�섮?�����ڍ��=}���j�C"7OE��U.Q�[7�����o�Ǌ������ano"OD�ƺj2)v�Ec������n9ȏc���Ƈ%7DCӷ��H�K<܂������U����r8yg�2�`���5$.7�Q�(��c�ח�T���E�Z���Vn��KVQ���"Y��)�������9�6�&��Q�~�]�-Yd���������wR֎�R{i���l&u}hl[GG�|���+ODn��7Km�t9Pj�����PS�pJ��1�rQ �@����#BUK���H�+�m�g$5.�,�C~޾�%QO�xU�z�ߴ��s3r=��1쵣���3�2r�E|���&�k���f/Q�d��,<���)��p/P��8G�����<����Ǽm�Y>���V9�p}�m�L�ԁ�ש�e�PG��,|W%ۓ�d_�Rcg��}`G�~��Y�2C�Z`Ic7|�B�Ww��(E���}O���x�S �����=�_��@�L��t��o!�|�W�􏈩��9����^cϙNw�5��Ѻ��bP��)9�8GJ&�s����dQDМ[��J�VZ�j]���T�t��_�ġc󝦤���A��fr
juB�uv`n�5#ӹU�&��,��Dl,��O����M��o!d~��ۉe-a�
��D�ѷ����n��E�0nt�@���.�&q��	,��%��o^ �q
�r���7D}���D�3\�����-A��Ll��)+9�֎�u.5x<V���dJH�Bۅ	YҜ�Q�Xi���(��?���E��G��oJw�n<Z�~'�ar�S�g�o�#V(	�T��GNӪ�� i�� ��@6ӎ�C�>�;�k���j� _<�=�����ꀟ�E�G���}ڼ�N�������Q�Ԉ�������o�~N�S�z���,>��e{X�J:���D�bK~*��V�d�%��S��@�W8����V�)]%=P� �R>�a$l:;�9���^���I~�lKt�$_�*�< �Z�8��(w�3F�l�I٬_��Y�GO��~bVH�{]�D��Ӽ�[Um}bK������P>���"���l\�v�燐D����+���l"K������<�W�T>@�S�r$ߏ���߷Y<�մ�A2��,	�߿K^M�;�@� =ӳ<<Ϯ��2�w�:�5&��b@W�Z89��Od�
h�,�$��T�I0a�s{g��bVgs����uq�uK�DS(�*��p�q���2��a���3��4���B�y�5�^���H�j�������`��H��{x��K{��J�g2,�65Ƈ"�+�x�۝Q��:�i2f���\��&Kr�t�S�#�J1�Қ���gye	��8�#�V��E�[j�)�Ggg�J.�ߋBk�vf� @Rj��,��绲��$�v�|�t�)��*%Q�T`��ݸ�y�D�m��Z�_쏸��E4�S>2�.��Ya:KyM-�� � ��ۚ�pG5|N��OA�����U�7��n�Y��z7.Y�zֹ؇G�����j/K��n�W���,*�;x��{M��8���٫�s��z�I��Wo�3�n�Q�f(���:�I�p��/�G�]_z;��&(6c�gN��Q�Ԕ����}I�V�8�k��HG�����E���3���0U�l� \�u�d?�����Ս�6��]�tgY�2 ��&r�߫4Ja�$vd<�{s�8�&s��1h'��}\G�_��G�vG1�H	�(>�$z��(U����W/ 67W���BԜ\��&����N��T��Z�$I������p6��o{o�cǬ*{oZ���֬��h��X����Z�RB�L5T�lQ���M��{����O���s�sߟ��9w8(�{���P�pw�[w�M^��䋧e�oR�aA������,Q���f2�f)���@t�⎱����"�/��#�b�3pԟ�{C[v����So��)$�%4���$˂�E��b���W��`��	z�@������� �q?ñ֘�_�԰�&"��x>?q���7�C��41B!�{3�G�F���ѩ�%N�s�L�{I9ӣ�y`ݒ��ׯ_�e�T>�b0=�Y�S��,�	Fo5��?�� +%�p�#��}OB��n��Bo��q�}oM	
��X��hIE<���%���z�iBG���o��|���BMCH�J���?*���{����_��OR�ݿw�yD!y���f��ъI0�=h�Oht;�8�g@F����uB��G���4}hW�3M_��Z�c�巘�=�`��^�e�����FJ��Ӛ�b��~o�ka%.�+�00y4ҴNj\��Q��A��,�jhh� Ү̊�����#M�v�fB;?2�Ez�bd�5�v�d|iM��G����eK�%$!bOm��^(v��������g��!���-}�Z'_W핓�R֔|�kbGI��0��9Ͼ9(d{�L��}��H�Gn�ݻ6���{G%�P=8�q�i�+����Ņ$�8}�w�A?�z�f`���;�|����ј�!X��u����Z��,q��@���K�L�3gxd$�qh=�I�G��@?e�/�)S::�چm�̅�V�I��SRW�p8F/�(��n����]�4����f�j����R<���DV`"/�t�M�l1ۘLso2�7l�#3����?mk7FU�*&��%_�y�=���?HbS����^��;�$�#�bq`�J�DE4a�����G&X��2B)qH����[�4J�:��	L��8�9���>���8�V]_i�G�GJ����Ŷ�����?�H|&qf�k�g"�z\�R�ˍg�2�Qc'��ƪ0�'��ր�2nN$164�]�$_R����lY��w�C�%�P�xβ26H\����i�}+���
���T�E������3bir�/�� �����?ݡe ���Ʈ'��fp����o?6ʑ)m��֧D��׆@@ù_q!INj��b7>�����LH�/�Y����$�_�&3����F[=-e���r��c�H�f^����}�Z�;�`�v�'�m6������G,��L�ms�)��ms��` Cq��
)b����)//V���4��_5F���%H�س�����Q���!H#�{��zy@��Q�G�j�hC&�N~1c{�D�
�뻯L�����5���:��K�����Qx����%>�\�7�r�6)�C� I�)aM%WQ�y�0����U�8n}4w?n.��\����u'�Rg́ذ�p9�����6����Q'�#�X�e��O�6U�ǉ�"̪~(eUl��Ї�'�'
?��w���L{����/[����˛e��*j���p��t��܃22�,��X2�5�H�x�w��32�Z%v!uhvR� l�����߮ͷ�ܩh]����|�?0;"���cD�;v�֌e�����X��X&�������y>�r�\��w�$\d� ���"��y�������tPkQn������,>嫳��j�]��D���b���+&tY�dŦ|*��<K�
I����rU�,�VV�o��t,�/v(HL� ��)���"�	-aY4�y=۫i92Z7�":~��M��6B�����ٛ"sh��-��/I�Z��Q۶@fX"RZV�y^Z�w�;��T��u��9K~up��Ǻe�=������!HB��e�m	�(�tyIw�Ѷ�A鸦��ǽ���{����x�K�]o�LЊ-�W�WL�=EN��)�6����w�):^*���%|���&�l�[�ܠBE����0.��gj�!��;{���Ꮐ��~#F�B�~�+y�nҚ�Q��R"���2�V���H3h�*����P�O�n0 B��b�P���^�����oM�/+w��l�I0��@��y��ek��#5d9<���Th{O�ZRmMM] ���}[����\��3i?���}Rh�z^�=:(6�v�*���L��L�pk;E��煮!#�W*��b�Ph�yn;5bQ�uЈC��_�w�� Ս�@o�6�u�	Qi ]��)���m֟��UUTJR����g��-�HF�(c�˄�-_�._ZZ"f�tEZ���\E��3F�6��)}��sZ=3qiG')�h� ���̥�i�����rޖ�QμI��{_�Ao��Ի��ć2�/���2�3vl���{w��h
�&5y��&52(kp�����*lPQ7K�V+��Vp���1~d�'Zd���|+t��a�SG�h�a_�SJ�V��pK{ ߷�N��m�5\��[�����a��_�(�춽Yf��+���6}�zrݨ[VMЍnuw������g�3���N�G&�1�4��lZ��e�M��o�z����u�Z#:9usK�%�	0�7ܹg����c//6�B@9o����%JJG�A�M���)��='U�q��~�jqTc}%�.ˢ8p2e6��ͦ*'�'�`Hw��'�m8�I_k��~Gm:չb�xK�~l����x�i��t��:�мt�Z�i�!��� ��&��G�џ�Z����ė��[Vܵ��kקu����
�t��B��Ovx;Z��2?)�O��ӿ�_z�@~8�(t�@c�4�G���k{  �ԏB/F�M.f�ڨ>&���vх0�
���e��\�(t��� O5������- 䵓�2�oS���Ĭ�75X�d��-=&�2���a�h$�w���6߽���)��j
ЁV�k�1ڦ9�s��Ɇ2����LV��VǲV�BkZ�?HI�ո�M-�N�*<ك{�����3���!)i��Y�aY+{T��a}��X����e�4^��O�`vm	�h�<�c�]���q�Q�L���##Rmɿ�''aE�b���=��˄X���l�Mt��-�>���	5�)��� C	��5�N~|eN�7ɺ;)���㤸T�A9S�LD��X��_�@��%-����j�v`z��Ԙ�FnsN?Y'�9H�Xh(�}㲅�������U��7��ڎ�kM��{�w��Pd�������]�J��ljIC�4���A݁�M�$_�$���J�S��>D#��/�-G�@"���J[�32{~9�2�������D�4|��L"�������g�
H����UM�* �C�������a�v�BƖ@Js2��h�H�w��9��"aeQB�E�9�M?i��4�����M�Ѻl9��t�?~ta��ˡ�U����ϑO
h�!�,Ȉ�%�t�J�i�5�nLѹ��S�k���f�؜԰��,�G�rQK��-\�q� Z�w���Ǔr��%Zr�C�s���+�"Ɖ��	y�<� �%"k��/5���+��;��t:��:9��;;H��@�EA�ܳ1|�`,�����lyu�@{��x���'WG+�����*�4���^���ՄfQ&y��F�߼Y�8�{�����"��FyS��iʌW|��@�d�WP�b��/$�|�ǭ$�����gf���Q|\o��3[WM�6�*���ۦ��ڏ�f#ꮸL���4�򁸼Xe�AfZ��a�Ǻ��y?ڑ��h��;f%���uT��#Y�4�Z��"���y�z*l���a�� i��CAĩոP������1��-\ԪOc�T)F>/�����67�7��O��ː�XoJe4%4c�˱��k8I|�!�.Y$(�b��M��������Y�_\'S#�hn8�q�r���|W
�nB�w%0}R��uc�7w��oU@^�k���D0[��{��=R�����JYLd��g�6��O����\$>FRC�m5e��"�%�Q��/.�$6���)H��e�<�>SV�/�q����݋�ۏ��w����d#Ť/�\�m�h? .S�Uz[S��oqflۏ�P�kn���ނЙ�n"�L���1Q�O��{��y��gfߑk��@�?���F�(�F��ȕ>l��(+*�x���.lp���JF�7�6���	֞���A��Q���
L����K�'2k�v����2��f*!r�KEST�6#�ZUOc�L�s�i��N���#S:f�/���s����J�I�N�p�lg\l ��� �{y����Y\d���~��%��4M�s�&'#>�?��b��Ĥ����?:�Z�I��:���dTU�k���Á��*
�ʎ�Δ��6��+�z1���5KS�e�q�R�&C>i\�h^�`ܪu^�z>I���,3���u&�)c)�S��a�g�&E �rS��=^8˥IN-gA5W�ހ��j]���60��y�����M�+PVߠ3�bV��j�x�ƥ_�a�esS��Vv�R�����񢑳'ZN3��ċ�e�'5Kj$7�;��q�G��/Q��|z3N���-�.�oV��$vu�e|[���kH�`(3�@$A��C$�<t�0IY�=K������j~t����{ll��Bj0�+�>�mIG�fd�;�Yi�D4Ͽގ7�=����UM��yzot�T}��k%��XK�}�B�/��(�6յ�&��|�	b�R��������Di_��=5*D�r���	q�_��1}�>�#�5ʧam��M_붙#Bm\�_"�͚����ݮcz�-@���j`�}���f��
v!���+3!7��*.8��.�������s�	|��X�^b��_��ۿKԋ�Ѡ]�q�R��5Ň�8o�)L+� ��_?�ļ�4�9�)� �im�z'�A�������l@��x0���})!�7�x�ҹ����{vF~�@��J�-��o�:�	�u�����)}Av]�g4h׏��wkJ27�Ƈm-�ޣk3�&rziT��
�K�,
D��w�o����M �YW�$t_E��YW���a�y���S����yU��� �<~n��ԫ�Vݹs^��F��k��V�c�ɨ�3�h5������w.�|1�cr{DN'�B��k~��P�MOl�l$����]ޠ�v)�ףE���p?���پ]ґ��T���y17���DX�Q���3�N�����.-���!P�Z�M��3K�we�6��nv���V	��adBCS�����w^�lpu$� ���d<}
+ºN~y�
��4��U'!|��+�����������xU̶L��`n�lb;6]Z���,;�<*]�Bq��b)=�+~��˖�
���YN���oJ�j�E���Ϸ�˔�
�';$.}�`�<�^X����0e�++'H�y�q�(7�g�lD�i����7�M��W&ձ�"�r��e�^4�|>&��Z���}���	�pw�?����^�+�;�ݜo]����JG����r��UB��hߑO����$�**xC���2ۉ���<vd�E���Qr�=�xW�}���e�F&�N!}F�l��YW��~B@��]HIsy�f�@�p����Q������|,�=�<�o�6�K�{]E�������B1W�O�b�f�R��rV�=ʭ�/kw���3b�F���I�~��}�>f|yL��V��JRI+*�>�S��C���#(=6*�p�~�钍( �wuŋBi�U�D5kY��i
(�z�e}���?��s���^�n����d�Z��N3*5�z[3_f�����&�b�Ջþ�0O���,�*��C��/g�����,Y�&�⫛/�4UΒ��p�`^��pd]���=�8y/���N���������u�Az�ĝ��!$1��E�#��ۈP��(ji޿�"�Bx�ڼ�9:�b���Dy���@���� X���g_*k�d>|����t�.k��ڹf�I�ʨma)<���S��V�s�@፳�Υ쉽�<�y7�p�sh����.��;��꿙7�;��F'������Q���9�i�3��	�zn2hhE�$1��Y�V���p��n=�^�h	yzg�v�;���ZP0�T�ۥŖ�Zd���~�����}��F�P�����򽍔�:7t�8���|g^U)+	�5Lxn']��ƿ��\3*W��^�C� �1��yV���s�yo[%~�ʝ\+��;�>��P���Oj�2Э��c^3�j�$Aj�~�@�@�j(E|���r[k�P�t$E���ǝ� Ȁ_�j�8��+�PW1�f5}�&j�����Vؔ׆y��{���L5��4��8�M6��r�a�}�g�r��:�/k��17�[��U�x����D�3΅���$�} �	�iT� ���+��'å&���D5��"����6�m\s<�Eq�m�t����0J]I�1����@�@���~�����|���y�����a�ۅr��>�ä���	�>�%�4��2%�7-ح>��f�T =�^F����+���_����J9߽ڳpH���~��OO2<�q���j�����G`2�[��eUY��p���}���!�-��x!d���2I�A����V���h�.�PH����[�L�g51D�v��\���tZo�Gɨ�w�PϚm��x>Y$��ߢ��d��p�u��;���۠[��bs��\�7L����sWT������*��pUP`v=3|�#)R�{C�E�Ϗ<L㤳I�)g�u�u{��$h3\���!�,Eh|�w$n{$m����Y��;���VK���p��G<U�f��{�|]�s"�_��t%��=���u�ha���U����H��=�l��9�����O���Ϟ�I�ްN����5z�����K`l�7)�Ǵx�s\��?vb��ci���Mc.Nv	ޘ$6.Q�7�����@.�_U�ӫQj7�H��	
J�\��y4���*k��ߋK]J�r_�-��ǾBHS����/�	�߆���ws�0�J$�����=����f�RoN���Ŷ�,�ڣ�x~��M��1G���Ɇ{�I
��uQ��Mm�s�lig�������0uu�Q�=��N'@d�x��T7�_th���#\r���n(U���~�`Ùfd�o�DA̞�zZ�&5b.Wo�,�L3"K0���{ט(+ȋ��|y��ݎ:L�-���.�<�q����6o�����R�d�,hs-����>#�O>���=1e�sItk-UgH#�^0�xY�/�+}v Ͼ?�m�y)���(V������xp��s����J�$�r���XY!���\_��j�v6�L-���06�BR�HF�$	4�di��ށ����?�i�[Ul��.��&h�+�{��-v���Q���=��e���y��mօ�}qT�H4�P"��������ʃf^�.2���{�!�T��5����ӣ͙U!�G�,EQ&�`T��Ȟ���y5\��j����G�0O��|��hu
�����=b�e��c���I7��k�9E�eB<ǉ�lII����d^�޺=*Rh�Q���6R3�P5IFa��k��g\�˞��2��h�>t������$&s���}ZK���/�)R%�6���o�e�D~��j3P��Znt��ܦ4�]�Zf32�pq�
��iq&���`"��Ƿ���N�����|�}����<�Bm�)"=&��U�I��b�י�]l�j)��l����O�\���;;;dfG�-kC-@�<��gCͩu#��INd�i#��Ա�-=�bN��vn�4o<//�4�O��~���_��K����70�v��v����-�-^/�M4!�i���#2"�D#2��u���$l����ߣ<�P�W�^-s��� ���U�9	�׮Գ�Ѐ	[�a��A�$����	e�6�{���N-�O�l�IC��_�}Y��\
���дs�VWL3�r�1�w8vLy��?hW渄﹖���s�*|\+c���o?�Q��2���y׳v�<����d�W{g'��ң�s�)���t�33\A�S��5:�}`�jF�6��4��0ae	�֒���J�9�i�����.A�.,]^�M,*M�rD�Ho��������d4���=�����2�$Ԍa�9��]�����{�������"a��o����/� ��e�iTڜ��r�~�H�xt2��~���z��oۿ�+����vU�ϖ���<=͕��5�h�]Q:������,�So��߇�2���4���faD ��#YX2�\L������q�W%"�Ҳm/2k!z�q��^��/������k3B�TI$d7m����&��N*��{]��<*6��-�"��iX�dg���~�4��^�
��-��.&��Œ�wÝe\N;{l�!�+��`,}��S�QxU�j{J��iȐ���x�5m=�)g��J�(���\����΋�޼�:�w_^�j^��u��ǽ���d�БV������]�?V�M£�]�"G�#EEW�Ԅ�� jɜ͎��W�)�`{�pS�{q�2�F�R�b��lp�|�>qW%Q֤?�&�4?�VdR����;:�X-꘎�9W|՞�3�����q��_�P��q���\�[/�턜�����ze�~�����4A�<��vf�(-��E�NC�2�3��0L������Qg�$��Z}
��۞�ƥ�;��YY�w<�Yd�)�j[U�W��G�_����M�ǯ�t,!>a��LC[��f`��e�ΙsyοG
��2Z�~m'4�ex�!Vn��)0=��ش�3��Ϸ��I�U74]y���־ȫd�q��.W��Q����������JnJ��e�P9�*�R��:�=�om����c�ۻc�EV������߿ɸ��w��8ؖ,q��������� d�w��|�h�,D�X����q}��인-U��I�[00�ˣU@[{��R��%ys���Sy�q��H�r��q�:�R��K���Y�����`^�	_��I8�U�n��]l���Q��ߎ��V����|����ND�E���否'��î���]�ce\�I���c}����O =94�Z�Јrz��G��TV��b��o�#kH����l@���H��0��0�|�fz��5e����o����lVi4��@Vl�4i���4�h�*��qFǐy�_ه�a攦��ai���4���	���G}<�K��[�m���9K�$����6hI�*������ݛ�ͫ����0����6��,7א?v�q��SOOƆ2,0F>j��4Ԕi;��V/0r�=+㰅�s�S2{]%�;W�9-��-mI���Zï��V����_�^0�}�j�Ɔ� l���{h�hYD9�N��ơ'��f�!���X�<KX���H�b����K���Q@?!�zMs� �ӏ�g�w�����]�:[��3sxu�K쎣���m���cp��x�[ި���YβMmk7���Td��N`>��w���� �m�/V��i�ϴb
�A氛�7��O�@M�����cUqs�{K��c/�\��}�`������<���	��&	z巒��	jDB�i��]�ė"���]��;Pqa�8�~�����/HZ55Ī��Dr�Q���Q�$�Q���
�����H�~�����f��W��DB6�ms��T��,U�ǟ��>�MR4B3>�Bg�e肁|��	F{z+g ���B�,?焞4{kh<���3gK�Mصˇ��ҕy��D��C��~�,���~T���ayՈ�^�������_ܦ^u~�^�B�t�����Z�ޮB�x���,\'��cO�C�a���U�\O+�g�t��>�u��b��Հ�3�S�n�􎘟_~gH�?K�b*�K��n��rf=<8)��3i�F8�wAg��\�φ�D�TU]sz.�͞4W����C9Q�0������s=&2��_B�_}�}Jʰ��ݠ	_q)4��Ű�)}ڊ�āLRb����C<��*w�=os�Sr J�	�1�f������Z""w��qqS��Y�C�;�Tx&j��i��`�;�Ps�[#}a�w2�fZ��6NŌےۃݽ)��.&B�uZ��t0��#�8���E�7�G^�V�p�\�f$Hգ��o��X�g�7��G�P%�M�d|�u�BH�/f�*%i����Ɉ>F�(���=�z�RZ�c���C�C�o$�J��D�A �s�3>�&"-�a N��l�uK񱚺���* �AƘ��g� �7�6؀hsV,v���XXpmQhH��P��H�b���N���e���Y�Zv��#�α;��j��!���h4:�e���C���m�[KI+�䓡��N�!��⛺���_̒��V)B5:O�(�Ռ�sN�r6e+SL8x�M�y^��p��n��~��q��ɼpw�a{�!c���]iq"p�>D������R��ץ��[�Ɛ�$}�
��\	�/�� J�Y��gwmj�j��`��&�\!���݆�d���K�9 �<�ڦ��'m(#m[8(+�,�1m��\3��8������-Ҵ�V�`^A^�qV���X�!�@s	�$��5k%E�������C��w��t���Ě����=^��?�M�� ����e;����+�>l��������D��l\!�D��� Y�"�5�ǭ�Q(�γ��!��Q �֧%�j���zUK: �9N*��b_�k�9(<��_#���E-���A|^@������(n���;$��ICo�}����X������PRSs*��V�JF�k�+�¹hl��\���s�����^�O�Ӝ�B��pwī(uS��&�ԛWW��|u��AssE%�ֽaȾ@�We��Y[�$���_��R�����Sv#�X}�͙H��ݟ� �W�ӡz�<�k�X�sw���t��gF�O�#���@*�Wo_��5����Rj�?a��x�Ў|�ޥRM�y��~wJ:j��ȜI% I�1h�te�
b1���[�u�� ��F�ZR�����&�;��������i���FS�tto���������_iR��|-�Q���z���E��i�2<�3;�%��B�i�}
�["Jp�V��% y�
�j�����S��Rg�b�wm[p�8� z�9\���U��ռ�U��ﺛr��7�ݱ%�=]#.�ܡ��|nо��{ׁv�=�K�V��G�dE�C*C5�]��2��G��������cR�KI*�o�&���4.d��T&v����	z����s���m f`��@��sH�Gb��4��i��� ��һTI����6:��D2fW�,Ѣ!�©k�N�� �&�Dz�y27-T;i��Z��p�jM�Ik�z8?�l��J�=�*��T$�U�t���qI���s��銗�Yjdc���%q7e/��SJ��4�~<�lgcV6�s�L�nHj?���a�d�hM��LGk����]v̏��,�ľ�f;n� W���E�3�|p�[1�<���j���s`�yo�����`-A�+¬���d�O���1<%��Y�(W�xu��eW0Yi�\�ݷn0�� �@j����5�4{�-��?������O>wA�B>�KP�m}�����*#��+���2	T?�_�R%��/�����������q���ߕU�\�ĭ�Y��nXW!������цL�J��ҁ3�^��Ɯنtv���-{�9��ȴ��Y�<[�Zz�ӣ�۸����M.�?a<Q�JM����5%kkmc�=Z�)��:�C����Lq�O�ږ���Z�4n���Jx��4�>�'��!+�٬$�u|�T`l,��EӬ_Ű����}k5ۀ��*��-Ư�B��#D)�CԔ�;{�g���3۠76�n���xr"k�PB,W�CpVE�t����	�~ේ:��3`u����Vy��`!���;g����Y�J7
�[�ɤm���c
z�so��η��We���1o��#"#�����j˛ui��Z�t���J[�F��y>c8q��ףG7�q'7�G�����8�^�-�l�p�B�V�ۿ���?����[c��(��+��H�m"���e��y��S��9ID�W+����JE�`{F(\�m� �!���-��?*<�_H����ǦIݯ��aH#�dȏ�;F|'O����r�Tkx�����zj�u;�,|D͐�bf�u��2�������r@�&E>�s�ڄ!z7�����,�=K���+-���}>������Ĕ�Y��˱���wH������d�,RiGS�璿}R��o��ѻ�!���������_�N:{ӽ��q��ζ�+O�K�yVԠVa�kC�uf����W�CǪ�����J[�n�x��l�q���l�C�M�g޷^�Y�ӗ��C*j$.H�	�$8Hol�.ӄ3�'6hx�<��쵾�e�q�F)ZBJ��q��u�f�Z �''�Ğ���W�E��O���B,���%�@��M��}�)�a�/���£�+.�'m�NX�?Y-�w�V�ȗ8P��ˀ���V�QJ	�B���t��{X��5Ǟ��ǯllP���w�.B�� �ߧϝ�Po}����+q�T�w��f�$�Y��0`&US�hѿ���f�C̓�%n�k��_`����l���]��
����e�Jl&�M2�����B)C�$��ش�5�.�F]I�X]I�V��@uK�g������+�0�e��UZ�5K�c�l�I��v�?atcΟ�i�9S߾;Щ�3���6�lhB���L����|�5�4�\���1����	�{-��{7b�R��Z"@@h(7�jY�����o��A�7�&�sPђ�7XG��E�((�їz���Yt� ���<}	2u���%H/��@˝�|f��9�d�S�iL-W���x�x���C4X�1✞�k�k�8�2Ӟ��;��7��V?�$�@ښb��yo8_R
�!M]�d2�����ŲM�X`#�8���N+����эё:p� �4Bw��<�e��s�|�o��z���O����!��ъ0
�]�{�c�+�m���S?�
�P��b��H��6�T��ZȝQ!�"�Y�B�Ș-u�m�I��|�}s�#k�^�:���Pd�d�zUV��6Ӻx!l�!�aF�w\�x�͈�WѬ���l�A0��̀���i�	!'��P��E1��K !"ʏ^
�}:�d�
�x�AY���j-�U���(�U�|��U��l��i\�w��R�R� �WW��D��5�_��Q��w�$T�KK�l�Z�C ɤ�J��S�f�dKo��{�7��g},��󦱯�|v	LDV3����}�w�9�z5�l�NEߌ;�{��t�����|�5n2��H+��[�ĕ&�]~�I$V�~��?̉�3'�
���W��d�Dir
{Ba������������`p��B����;�B [�0�)�5K�=yp??S��(�]���S�Xu PhQ��T�)Y�,���-�\���y��q�{�^�Rw<�6#���J�ZDxl�Ba�w��H��7�)e1�_���Q���wc~M���*�����azGGo���7ٿ�啾s��_1��'�ZL���BD�Z�K\��-rm�H
��4_5���������"�����^���3���7g����5~j��,z� ���ZM����Qd��֪�'A��Nt��f8�]����l�=���Ji�/kb�#,s�|p?Į���¢��W�B
�D��.B��L�{B��ע�'$q}w����P�%�����;ݧtW�G��y�`_������T`��jWՈ�(��z���m��z��8�x�zF?��Ӂ�Rݏ�X#�C��n~�|>#: ޔ�-�#�.�w�Э�&��>x���v���CWx
���Y����ZH<��^�������˺k�k�d8
P%i�L]:��L,\��u�I�D_-���|�#d�����4?0�柳��n(_
Hg⧶n��֬�$��qI�z�J���Υl�ĪS�R�T��!і�.N�Hl��Sj� �����[�ä�.G���G��|?���}��?=�lH�QRP�!��<*If��7?'[[��Y"����M.t�GE4�j���V������/ْ��3�4F�-/퐚�=��~���p�\i�>o8�1�2R�-���C[�Xqi�u��Ɲ�i8BSS��4��<3���`ذ^��m�͗Z��NkѨ���|p����-*p�GcAi9+�q?���˨��Ӥ.���9o�UBR�ɋ�S���C�߀�I(t����r�I�h�����[�4o��
�"���9� ����KI�ΈcƁ�ń�7دƾ�2k�P'�1��1�^�[��w��l��$�QQ��e�sw�6��)�9�ct�Tb��z�T�+;e#o5��kGH���~4Rxz~s����M���œ��5�Em=�9�`{ݼ7�Yu�^qF��h0��^B:�#h��������z9Ay"��?�ΐk$li��E�倨�O�8���s����XB��b(!Bsfy B�a�da����=Q��k���ώ[="�@gy����K��t-��b�`,�NPx�ɴ��T��ɭ>]~Q�w쓹���ms�St��#mu�C��i?�d���}�% }� ��hOW�'�
i��w� ǚh�>�&��Cį�P%��K~x���k�jd5��S�ӣ�K�����'\������(K�v��3#�B�;;GT�nPu+-���g,+�����dca��?�����5Ki��3�H��!�i�F_��L���y��Y��� *^/_
<�vz�&y#��{P��M�%B����s�������}�R�Y:?z��\As'�	�A����ȹY�JG��X�ը���������h����ƝjƆ���1Gk�e��G����g�>���戧�mV��2cܥ0��_�6�����q�u�+&�l�5���5��8��S`�LE�C(���#�:�K�L1�vx�0�����Q��B��kˤ,A�Ɲ{Ҷͫk�� �B?7cu�)�/JO�ܺ��������������0�1��9�"�6J��M�P:>���=�M.}�]�D"�Q���J�>����7ݬ��JS�tȋ�Д��?ӷ~h���oEn�y�G�	��#�x6c`��2�Q����(7��FU �� �w�?a0I3��>�������6��9t���LTd(�\��;��Z��z4O�z����@+k3���JH�;jk�c:�qiß�������t���+v��酑��/�@?�%)p�N�}��ͤa9�5���BYLܯZ�}gD.�@��Z�e�����Z���+jB�ʘ�>z��R�i7%{�/�OI�c�Օ�$��VGS&>X���[�R#k�-<���UB�1��`�KrX�EKF2"Ԧ��*�c���/SX��ԻUb��ő�z�Q]0��dY��~.Aɛ�\n�P�����IeN���f�,�]g�����㵈�H�B,�x����!�"�݅�Zxy���o`�q�,T@���5$\�aX�F�
ߺ��@�H�b	�i[�_��`fϔ��<+�	��ם����0nj}��v��[ c��À����ިb\2h��!��w��,�K�!$�O(�m�<-$�����:Nd�H�Ϟ8J�@5���r]8p����T�.zy �jKW�w�I���s��d�}d �*��i�Z
Us-����*Y6~�L�c;��Ā@A����Y�ڢ���L% �������N��_���� HD���R��8T�@��`����=ݫ�)���R�6���e��fR��A2��L1c`�!T"v�{+V��w�3�ho�y�J�����6d��ny���~c�3����E�o�)����ѵs���~�� 		6�q���vyM܆�X1�ǹG�S��!I͐F�����8=40P�!m�(t���fΤ.6�A0"ꇔ������ұv��y[4�NX-N�ߑ�;�#�����j�����K^~c6��d�| Ԁ����ם����e&���~�g�2]��1���L3�4�1c��� _y���?/n���MӸC�	&-�JX�-uh�Z0��U���C�������U�iI31e�^	P�\b4/I��*sy�"x����O<>}�S9Mz���NySV� m��m��Ѱ�`�b�$�K��J& !�
�����&;|�<����K���K��5pP��&�MQ��3��筺���̜�-\ݕ���O�-��#S���Xz��*Q��+�:W̟���C����u�x���^f���B�	���f�8���C��v#��9�cԯDCV^N���sf���]h^���W
{.E���������M��hN+���łN��0��Ֆ{�Gy�z�Ty�ϦԠ�C,Vft-���	��� �L\��&ȔT�̯��oiS��b\�FJ�C�j[�Q4� ��,�W=aC$�s�Cn��t֮W
�_&�}���	9���CUA��`D�@�+ "%KIP�WK��.�V�ܜݢ�@^��LF~���� �U��
�T~�Q>�X��:6����{��	BQ4�l�M��Q��K��E��G�ښ;�&4F�5R�K��Ek��������I���������u��jם�P�b#�w�=�Q/٬�$ZZ�YUӔ�iw$�k�ܰM�}}�Nb�����A�( ��U��z�a�&*ȝP��VG:��0��-�/HŶ?~0��T�&+�\�����P�94z���"ꆏ?1V�w�l���Uٰ&T�Į}.�e��u#�!Rd�r=̾Ďd�
*����B5��z����-�2�u�4:��<T\���:��=�׽������7Q�n<������_�����X�i@��|1�٤_�v�;�l@�A���G��F�����h9��,!�A�����O�L#鐫���'�***+��E�:>��U�Y�;%n��V�pV�zi�c9�tJL�$:�@r0�t���Ɔ�ȯ�w�E��E���^J��̐�%|&��W}�0�5:d/EKp	�\�Q����c��4�"�E-��R$x��y��2� �7�y�WAZ�S�_��O�qf��Z�\`K�J���8�q5��%��>�'H,�������x��~p�e�yG�{�&�&��`	NF��XX�w�7��6=�/:ܔ��c1��+���������VH{��@B��$ܵ�.�G�_�[��s�Ч��u��U��*���}|ۭ����D�����H/*����%><,�U���^��a�Na%cII�t�D��(����C��-��Υ�~���~�m�鿾��UMXE���"#�:;�g��>�'���P�����[��ė�ٹ��8����8��߻�!.�v�A<$�=�h5JG��:���s?��&���%&������'nkϒ�y�����_�L��M�`���<Lm��4�q�i{櫛�|J��z��e����,ȶT���q��ݙ�x��=��r�\*r�)$6]U'�]a5�xIM
Eڐ�$(���M*����~����_U5��8E�o��&$���\�kG��A���hn�Yv;�����/$q�GLz˅�$|��:�� Q��K�}�*}E-����$~��<z����͑�페o}ͪ��gK����U�W��ʜ���;`��#�^����[2?�:W��e��z�$m>'�M��@ 6H�0t���r��u��p4��Y���/��d��W�{����}9ꮿ�;��Fɚ�`�/{�nYx���)�i;7��r����i"&�*�rJ/��9U	��B}u��;��4jT���8_x�/�����l��֖�_*�s�����e&��VI޼y����p,��:��?d{�Q��hm�CV����L9���y�l������ ���p=e��/P~�{�dT��ف���2���+w��긧ۜ��3B��h�E t��n��h��?UJ�ƞ�f�;���ߊd\rm�Jt�\�R}�%dP����78�]�mE��ؙ�ct�e�ߛ��8&�L0�B/@�`M��@d����#�~J�����ae�d�7��X���q׵?t�g�ݣ���!��&�F�[�0�i��Fx9b����~������\��7Iĩ�I��l%c�! �Ғ8��Z"����d؀��JU2�,`�#h�ϯȻz��{.	r�+�T\D��~�Z_'��B܌)$M7L�2/k�/��3��=|I`�z~']���Gbd�Ő)	���4� л��9$��eH�a�a6�O8�x7\�D�ʭ�{@�
���_S0��j�%��v.�i��[x���c��<r�	:��H#�@b���in��*�
���|T��Ё�m+�9M�Ț�(۶X@rI}�ç�s�F�T�w��!�`�J_Z��J:�Xi翡���˃)t�?*���<,�66&׊?�۾겆�ISL��w�Ǐ![�xdQwP���_�flP� �Ev�ֆ �ᅰ�G��F�>C##��X_���4�k��WeQ������D�>^���jw��Nߋ8u�|�/J佻"���-���}��+���=ܦ/���ߋ���9`����Ym�b?)?��?��U
��n�ğn�y��&��v~�x ���<�ϯ�-=�͗;�n�]��Y�����:l��{s=�̛��f��d���;S$���Ⱦe���wpċ�I�M�u���>.��y��~�N�H�0%�y�(`��z���N�v/�KyC��XOc�m�~_��Z�<���yx���Y������DD��L�?n�2�S��3��uz��֯E�-��x��ײk�BY�sBɜ>�&"���o���|�)� �������&v�ؤ�;�����K�R_���2G�h�W��:_o��f�ue�d��2Z܂�䇆��Y��5,ྚ���$W��z)XW�3c���G���!��j�����,�>��E�<н����D�z�,ߤm�������	���RO�ԥuJ�=حd/t�߉�U�8�c��)OǤ�����yj�1����i,��D(ǵ��b�r�J���(?O�%�����B�]nNg��8�q	�$IeI��A79���RI�P�oыQ��il�u��0|���C?��/����NU��r>G�}������>�+a����/�ca�o�����s&m��4H1	f�'�v&Q'���ػ)q7و@&/1�����zz�e:�vr��J��szĝ�)s�wl���)�ƨ}D�K#2qD��rf��}�Xy������Hd���-bE�YS�'�+�|
]!�7�gHoa�����[?��qc�ǔ����Ҩcʛ�����uؚ�VVWK��KfV`h^p�F ��K��p|ɁLr}>��-�L�Zߡ�w�fbΜ��W��RN���$��s��\U��O�޴w�`���G�(� "cg>B-_|���[S�Z��YqIq9�CI������]Il�&z���E����J����TT��m�VΗ/��%b46����ٰĳ,����o�����|�o�Ϳ���B��:������b\ ��Y�N���9���j���'��<�T�y� q���]��9��
�<�;�K�C+)�~4c�q)�!�}Qs��Kۻ�]��{E����%"��U/[˪�Y��k��"�+��.���y�hi���Q�x���x�y�(�cZ��slސP/u�l�4V��5j ��|ԥƭÑS|�k_ő�i�	�.lg�6�m�e8;)�{�F
Z�aB>��i�^w_�H����?G�O�/����{{�1�I��U~��[�L����%���f��T:�|���/'�v�@�V��h�Z&8���z[8�ɚa|����3(�4�\w����sK�_(�(����N=��e��������d�n���;�s�7S`��s���e6c���6�Fm��o��%�^�2h������3�:��	P�P��Q���CM\�F��֏�+͆M��&kP�A���]�]��3�e	'�Ts�ONm�{�/�ܺ�,�G��!�]&Y[Q�.V�����bVi�����Hk���6h~ku�2�Ps��p^��v;�ȍO:�}c8�o��Ox��ymR擰���h�<���~L5�]Z��?,J]���c�f�,��vXQ�V�%��ßĒ�k�|�Q�%�"��Ou�e�bP�������p�W�&�x���pʲ�(d���ģ�!A%��,OO���'e�Th��3��YF�\��o����`�O��6�E�G
�:(Р����݅r:��wzǪ6�Fߌ�?q�>��xV����ApE���F��Y��֜�$��]�iqc4�VZ�tt,͈��:b�s��^V:Ή��,�B�z��������.E)�G�P21�H������{݀�K��x7�V<�ˍ�n�#�gq���>�)b�K��3�|Pk-���M�'5t��й��]����/�J��Â�ў����f��x8u�6ϭ�8�Y�(����������ֲ����[?T%M�~ж��ꬠ�-Rj-{q���d�6x&#%�\�b7�.�T�s�;kMo?�� ��� &O�$��MPS��E���%�w��c�l��P_�/'ҝ�5ؘ�7yޚ[gvAE�!�y��+UG@��]��-geV5e~s��_���e5U��)�i���@�8Z�C�E=+�A����#���X��$���4�aň�lT��J*O{56������%>�Ё�h��ꆗiM��F��q��J���<^��J���ro����C,� ������t}n��f�m%<<_Lɍ�%���L'��݆6��"����#��*�]�ӣ��J��Z��h@�4���]�A�F��e�{3f�t��՗Bd�Z��T�,`��R�m�<�I�M�DSC�Ι�#�m�U���T?:$��Gp~�5#��1��(���_~]հ�@��Y�ig\��76t�|Iקr�B:����<��e9`�)$z?1�I��D�����?O�X�q�Is'j�SP��$��q�5UD#=*����3ЌX�i}!8���#126�����c��!s��>}6:S���j��ح����ݝ�̥X����н8g���wm���?Յ?q��2Y>yg�'-������@����o��*(�j.��B��kt�/�{�]8b�zس���P�P�]�Ӱ�8Ίx���e���ƟH�p�s��hQ�~r��{�I#��G&��s�nb�SP�L�8׼<x5R_
������GVQd�ޱG���i�@���
�={F���p�\��R�%�b��La�\v��tl���\o#z�?���*�9����q%��D�T24����M5%0vB�9���
=�����M���� #D0��U.�~��.t,��,�b"�䆋��yiO=ɤ�ϝ����|.b,G���,]�"p��O	9g�"�ɉ��%gb-5I����Ӏދ�ު
���\&j��H��4E��~��4�#9/�J�:���#fy�Fj��s�k�m��g�r�gU�ҋPo�T�l��-߃���6X,�U-#��J�u�yK��j;k K ˝Þ�S��J.�"suS����M��}T��&���"1�2/�a���.WnD��WH{Cp���G�3m��.'YΕ0)K�v�f�W��tN�(GSR��h�D�b��������Rh �pX_ovS��*7���ki�����&nD#$C'�j�$��YZԏ�aG$��(1�:�li����۲^�!���?u��x[Qbt��$;`Ω˗*Qn3|�3[�C�d��L���"�ӱ�Ub�s,�4��˼99�B9&�=�H�wJ�A�6ae�f��JM"tN��,�<9��/�}�b1�˵!��n�����p2�$��vYäAҩ(�Ƙ;�J���:r���1dޙ��\h�<W;F�ƴM���,Jj&�*7\|��%�����;nl����}A�����Ni��-H�i�S�����v����t��R�vS�7��0tI��&W��d?�A=�0P�4��Q�ݎ������ר��M�ʧ����{_�yhٮv8;)O���N���}�	�1gE�g/�����}~?�||��i�����g�-.&`~��EF�Â��Z����L���M�RV��B�(�dq��|����
AP.O��c	�̃�ɠ���¹��*:��B���[�j��9Bh#N��7����S�<�YB&�6��L�}	�j�����vױe?a>���@���}&�@�T��݆%��'�� v�ظ>zSkR0D�6� /m�˼c
aq�r~��|�u���$Gv�#���@/���l� ~6,�*'0��H�Q�-yPE�'tT/WOWJc�!��7�<\�5��U�7h�;�]��-�]��YM�V�p3½?�� �r�E/�g�02��cnz���0��\��Yz V�'�n��j�TH$p�Z��*U#�|�S"W#T�<}��
�����mY}Q��4<řlpI�TP��ڝ2rNC�^sΉS��OC�iyP��S���"2�Z��^�l��,�3�K�d�q˺�X���uR`�J���L��jY[@X��t/E�v�f0�����~
7�,ӣ��e�f�{��O-QƳ���V#�iENV;����Xr�b���`{9'lÇZ�6y:!���@q�ex�w�RPφ����9��KS�C�ޡj�AmD���)��������\]D#�^�K��[�����{��Hj�h��BwƗvI��K�����2�1cL�⿓��gC�H/�$����v�=����;0�Tm�]�>ӝQsr1��M���#����g� _-�QZ�-�4����d�n8��Rv�a�~��0�E�NW���������,3Eƚ�4�KU���n����o���L!0�is v��;�]��=&J[��\I�"�Nz���Ӈn��A[�&�$��դ��4���
�����10;+L�@|,���{��چ/C��D�bfb��]2�tK�"ߙ'�_�ӟ��H�/�E�#��c�V����?{'�z{ڻ:��Ӄ��\@��1f�w�R�;~��=���[@�H�M�vw����a�s��5!������p
]������?k£����@�������j8k�>]t��o�ˌ�68S- ��f$DC�����^��A�&[ZM���SrȂ��p8��҇����*��0�O�ݵ}��e�&8�����'J{��"2�8pb�:u�{�fܘs�M���U��p
w�VN�����ui�B�����;r;H�$m1�k�ㅗ�0_� y:-�/�N�p�b��]���M�������"�,�;�j�l��&�#�y���Ű)$^�8���7���Ț�qD��e����+�sn�L�]J����,=~�%�n(�z ��g)�<Ҥ�Ԡɚ��k��[�0�ӅZ#����-�@�Y?��������"���������@��/A��P��v@�;�t�Y@]����LWnM+��f����)���@:_�3'-e�hS�g��� ɝԓ�	�DͰC�Wc��\d�K�����s�مm���aj�W5p���8�Yp*�uP׎{�5�����p?�&h��nw2+���_���u�_о�s�Y��@�<3]t����ں��$iS�0�` 	�Ro��K�U�����Xu�Rw٢>0��aI| w�ʛ=	�W��醢]��.҅���}����>��EQ�_ۜv����ZmC�WS[2|�4GF�Ei�����ʁ:T����S�'Z��5m� W�둝�T��>v�-,���x���5�/�&�9�w������wn�$���$��@��Y�����<����z��8߅����҃�	�Dd�C����,Y�+��o&��ʆ[�~0�2��6Y��/Z7��}[{进{Wk���������>�iX��&ߢݧ��M�ί�+��_���IO#dC�XSH��Y��n�`�A��蚇��)�������^z��1�e����h���tJu9�J�����$!�K֨�~ip�{L�ĶK�{|�p��I��� �g.�!�9�ͩvx���oS�@���~�eJ�'7�Z��h��-�9�@ߌ
	�$YT��D��K� �� S�"�t#Wv�s{�5g�"���|��BW̚/=�>�%\B�-�^Q%d�H��.�Ϝ:� Gi���^��.Y�B�?��r�y��(�=ײ����e�4�z�%��1R�O_�Ļ�a���p�}�� �m8�1��0��h�� �$�l�]�~Z�st�q���鈀���Ǥ����C�i2S��ۄ�����
�?"���e\Jю��SJڌ�.m|q��u"(��d�OND9O�q��t���ѓl`�o�MZJ9��f��&]n��~�Pb�ߤ4M���3J��@�=��ߞ�L��u�ĭ��W}I�����x]�9��%p�ɆlC}Ęm��W�&q�~i�H��K���;zt�]���󓒯�a5̵]�V�HS�@���9���	�j��WU��]Qה{q����a�t�V�,	Qi��a�����Yw�q�P�YR�q��K��%Q��$���W��>�H�����{z���yyw�=���kB�!%�����"}-!I���յ٢���J��Y��
���@/Rє��2v`" g��<,v?8�S�aqt��RY�h=�@�l_�mqq�"/x���t	��.JY4 ���W�&}���@1o��0т!�ܾ��&_���Q�wq,���z#5�S<�}��麏_��a��=��E�w;��gl���us6���:�/�e��a����L-3 �d��㿹��yf�;4��_i�N�%.i#s�W�K/C���4�����5\��3dK'�tA������ϵ��ǘ�Ԗ��R�������$��<�4�'E"Y]�����B�yR��'oE4���ۻ^�I�f�T��������Uޔ1ږ��P����>���������H�;d��,�4��Â �W��ƪ�!�~kx�Q�k�y�uq;c�v��M!E�e�Ò�C{K�A?S��:����P�q�o��!	u�Q�c E��"�����T*��yqu�H���D�������{cj˸�h%Q8����H�Z^�\��]�@˴�o��D���8��;�0���Ƿ�u *sl�妿Lu���W��j���F4��֌ ���r�2�?��T_�ր���Ȍ< 4�y������Ml\�1U�8Ym��uS�ɠ��w�pcf}"#<����R*}�Q
�Jr��bĲdkR�x�Ʉ�eɞ�]<^�\l��L�nM�`0�����_��� �l�v�fq���,l!8p�n�oU�J��9wր8��8
e�<�xr.m,K���vN��W�e||S��҇���F\4�??�J�ap7�8�!ԈV.6*�%Ã��2�f�|�n���V8oIIIȸ6����]z�ߐ����}"�9�	'ї�`�7_&@�u��ۡ��C�/�iqq(/��o� �۔�G�˷�X?��{��2*�z�j3�T�vV�Kr]�L����=Z�C�(R��Ƕ2��㢅����K#����9LF.?޲=~'qg��,As�6��O=�9�
�����M�-�+{{4�]�N}z�\�1�^�K�0����T(]���B(�s(F�����$L9m+��CK�(Bz_�PBl1'�3�A��土��N`�)��4�5�|?��XN�ڦ��]����̝�	��z��6tBd��@԰�z�)���m���=��N�o+�yf`�8����IMH�|��i�d�Z�6ƟD'�E�R�Hf�M�Sp[��}����r��:�@_�1�{ {\�?�}�lD�����.�Ѿ�~�.s;��j�� �r���x��7�B@�]�	�W�E0�­OQ@l+�A>��8yjڡzL^Μ@nuz�;?�l�=[�9ߧ�ݣ�&�pI��'x�v:���|o��H�Z �l�5p42~�r,=����Јo4�a{�|���]t�(�4�ym+�椓
��Ѧc)lK��}��ZT�=N�"F j׮i�7?u�=_�AOV���o��k�qu�׈K�������$y`�q<wQ���N|��zsK�l{��R�,y`
�#���t������	����8P�MT��[�W�j+�05�t�ePM4ń�xn,yv��~�G��6�dn��t|���蜞��0)nl���m��{�,�h��*wS7��Z��Z��?DJ���o�L֏(2��e���qH>�'�5�Ğ�Ti�E�U%%��-lm��LL��c�, �O6Ч���S��@�)0�8����2	�+�t,{�8;Y1P1��+>՞@�7��O�乥�c��Ij����J�
���\P�u�g��E�C��͢&��c�?|L���7z]��:��
_�N�tR�0U�~��V�5	�����sW��8W���4�m���E���®wO�q������-����٤�����\�f��$�u���		�X�����&�J�s#vu#t�d	T�9O:�nz���"��A�d��<���fc��rB^JfRg�k�H�
 �a|��m���,�EH)"������o+�} T�Wǁ�>����s7/ �mc��Zș��Q��Y�� SK�����Z�/&���ƻ�����!S0�[h"1�E�|�,m?�X�K�o�T�h���Kɦ��Ӹ!�e^����%(�Pa�h�~�tB�������L��܆)��/!�-��ȯN����zԨ�r��X������a��C��:���g��� n�.�8�z�6���!��hCub�+Gl�'pT�2���N�g~��х�߰7����yٔ{� ���AG>��~����duBO���6�r�t��aҋ�Y�$� ���N�#36��S�����XUK���	q=�H0�L�U��B=��T/U�5�Rh�e��X� V#�Y>�R֜qږ�0��lgo�@���\"�</�p�@m`�zj�-{?]b@�΅��e��>4��tKHK«0A��u%�l!�ާ�Hq��tA͏� i�l�4����O�E<YhM'c��N�j?�Vt"ȶ[
�	�MR������P�r.�	��i5��B`�~N�[6��!�W6���FXY¨��8l����~W8\��ѥ�]]�#�w��y�?���ٶ��M���d~����0���k���L��ih3v��7C���Ԙ,�I�`�B�Z�Gu�=��d��&�.��l��z���8�#�%���+��en:��&���7]%�J�!�;3Ƙ�ooKJ��:��;�ߌm��'o��R����\_���̴�q������:KP�p(74�X$#��@�����2ç��2�"Q5Uu6N3�
H�Nn⋇�����s����,u����7~��^�fI�9D���6E����(`O� SP������%V2v.����;�bYD<�bHy
X�=��c��c	HEGh��+���t댬,�<:{�
2���j�N�?�� h1�V���՘��$��Z1��K�(9�~s�!afMFn�G��Y����8�a�g��d��a���߄�s���{�o6�u�'��i�$�N 
X��h��bS��Gߜ
����^��i�+6 +���V~��������|�������Î�؞Z���v�Ql�u�ǣ�4����n�����S�sa3�0�=	f��vuJ��)86����=>~	��3w��-#7��_SQg����E<p烸x�����&c�Xi�.d���i|�@���a��#-��r�ܨ8Rm��ۮ�Bї�_�\��,�ww`_vI���a�%����")�\��	MHӆ�����Oq��
�=*����D��� Jl�p��0������7��ey��'�#�j���R!�x���������̍�x���˫{	��Q
o�SmQs�[_�2��V�����Fy�u�a���h���o�[�,�R���r�W�7�N�Y��E ��޹-�q��E^�M�h5~�aYD����|�xV,��MV=�br���l˪���/�-�_��r��Mw��{�&�K�x�J0-��1�7i�@�|W�� ��]'N��˥��ݧ���<N��h�9�_��������0j��׿5���h�-_�6_9Ҕ��Zb�ПܹO�8��XLe�z�~�ɃL���� ��f�+Wk���)o+X5}}���և��Azl�;*Ԓ~�j�L���`�j�F�@�/0P��2�i�C��;��9ɝ?���q�-�3�S�Ă9y��t�����ts/�����t3C��^��$($��s����� #�`7ޅ��2��f)���d�)Kl��?"�9& �#@�{���2��!��S%��v�tl�KD�J�N���s�@g��
Y��ҽP����7e��&mXG��R�=禥7͛�9w~n}��N���Rq�;�Rkp�?FI���9wv�I9�b�3Y*�"Ón�o��O����9���c`)2-�M\�}����7��/OD?NK�2�����7���@�����M���1�� �3�:O6mDk�s��Ь��g[H	�&`�����o̟_�V){;O*=?y��p��F�Gn�=�t$hM��Z�5��0x�nL��%{��f�n�/�Z�{x��'y����0<QY�0���	�̬Ysѫ���(UU:|w��X�Ѻ�%}�yH���i��g��H�C Th��D�b���T>:G�x|�ЂpS��4��k�ø����fOm������=���6pX�b�왟��ʠ��	X�3���Ibw�Z��MzgK����c���1VPI��t���5~�'ͩ �rQj�����oy���G���H�Y��t����ė�?��i��?��y��C���O,w���(0�¡���
E+��W?�G�/����|�q��r���i.�s�:ŵ�m!60��
Ѐt`����.X?OO�U�pX�=R�����,�s4�[x�8Et���j�toMӧ������*T���m�'���]]U���?qͮ>�u&��/i�Ep20�o���`	��r���G�ٟ�
;�|����x���`k.DL�b�a*I�l'�/;QY#�NG��^0�d�ir��W��s����f�ꞸytW>�x&M��Je"q=��_��y���K4p�*�S�ϛ���uZ C��1���/u'w]��ܗ2YH�����1�A����	O�������ҴG�Y+$[�j�<HzD}6�0�J�����3T�l$�Osմ��?V��Ī�g<�6`���,�9:�j�N����_�;ZܦV����R�OM���_�7uU���xW���8ދ'���/�z�~����e<�j���Zp�?���gi[ִ��.�H�[/�����K�W�e$bѥP�ٺ�bR�I���X�y��_��vTF��B���wAc�L�����h�E^��+�H��۝mYN����w�:s����K��>"ݬ� \]j���
/�}ǀ�L;�@0tn��2i��Kfьr]W`n�FJ)���,�L|g��O��%V�H��ᑃ�"�מ���. oH����s�ڣ%��g�M+w:�%�x����ub5�vsT�^"�&�>�Sz��/�����5`I�et�o�D�LT�1�jL�c�P��ylK~��Q�sI?�nm˪Vi9�x2D�ş���k���`�C�����w�}t�.2cUz�ù[�(b�K�^u��g�}��׮��~m�&W	=���N��=.�b�@%5e�&��QΒ ��V�tB?;<"ml�â��B�h�J����M(Y�C�n;�s�������06j���8������"�����򻒵����C��l]7�X��XG\��wx���W�vZ �4����HS��;��y���e�#��[Vnf�qz�$Ys�D%���z.��!�&o�|���d���DD=(6b���:鱄#~?��倰௾�1�g��	����	��V���<��'����}��惡��K3�NBe9, ���*2�D��c���R�xC��L��صS?��*ٱA�kdգT8sIC)X��C���}�֐����
�EM�>L셻����R�]���fZw1�d.:b�����a^�$v�odK[ L���y^�F>	�j3��o�����v!lf�� ������m��=���>�.���P.PH'������wv�S��F�r��
b:8�:�^@�):���9Z�r�Ubr�Kk�Cao�&w:Ȧ� �(�������Fߢ� I5� �0Մ�&��0LX�l��l]*>;t^xr~���L���_=��{�G����e�=����H4�p����y����~����0LqG'����hD�B��E1�"F�P�uZ|>���	�י�:2ߣ�2��=#WnѺ�Dv|~n-a�����]4A�����$X`�8�l+�mɏ�AU9_�����-��"C�/��u:��j2��,"R4˘}�z}���k�P�#�����^�⽎t�Z�g��=?lu�rcM�M��tJ+n*���@G�Qu�?�;8:f��/�������#�,Eb����SЁ]�p����ek��M�1�E�7(���]������/z�2����U��U�2���h�d�Κ��]�38'���L��jH��'.!!|�5[OA�H�WH��|�z����P�랐r�]d�D����uZ�w���Q��埩��!�y����}'��?�vJ��:۠�6������]�t�����<���t�uv�ɝ�e�F;�)��ʹ�J�'g�������7Nz��O衢����"E��3�CZR��T��O��~�zG4�)�^/�i��_^G?����_�>�k �c�_si,��:;;?�;�sc�>p%����|/�X�!r?q¦��UP�CzϏ&�UL(r�	�~�&�8�-���B�6�
ʥ���b�S��=��U�~'�?��T�ti,��#m��á�m�2F�ʩ�&�?F��ó����C�.vL��Z�k*�XK|%��^�g��Ɍ+S�H$=n�����`�I|��<�4g��t�,(��*���jw�끳�q�����ә�U�ѱ(��5����\z�ݳ��(7|db��:�e�Z�5�,�g^�:V6&.�%��VVփ�j�x��&-�|�x���E[Q�n�r�/�3�}�,]����Q�y��mx϶�-�~��Ӂ�Ǚ��e���ν�������wyWWW���Gq���1;�0����~'� ��c1CJ�?D9�ծBN����Oxoi�*1��q�PD�d�rX��>�r�	���r��x cՊ>.w!Р��Gr��E���;�������ЎٺTQRf�r�]���I���p��%V����[�SA�S �3�a�zP{g��7_���Q�v\jh�%��;�[l#o-�$a�9��A�;� ����JO��Bc�1
�ߡS�??	�yi�s}fs��L%�oA�\����5!�����6���M�D���q������d�[I �*����ۛ�6;��ކw�`Շ���c�ض�޼oU��O)��;YU#��?����nO���Vͨｱ��͟GV(�;�G�]:N���8�i��@�髍�G�*fe����5�/��.��~��l�uT��	vC����?����'��^&&�b=LG�O�-��ՔS��{�����K��S<�h6,��~��[S|�%J����̉�s3(�2a�#����WV��Qz@�����$]Y���w*@��v�3�Bǚr�|�z�,��M�%��=ܮ� ���r)�cq7��ro�fY@_6b�'��6G]%Ym�C�3�Vu��j>5��OV�ș�r70�˛��_)��H�mV֝~�3�?���d�%��ȓқ�h�ͼp�V� Ha� @�kP��%CK&H�\��E-��u�~��]n��ѝ�f�wp��^㛼��l ka��Vm?<�*,"9�����i��<w�9a���]�����c�&�(.�����}��BЧž4+�'S��q�����Zy򓟈��G����->�m-Nn]���0��}�к �5C��I��_o�T�)C&$6}v�{���N�t��m��q^��ތ�I��@3�Pg����+,�IAYI^Me��9�'���qw|���^�	��sR�Ҕ�����|�=7�W*4RB�y�<Q0B�6^�Gw�@�$m_%]���䷬d	�ʡ4�Ă^�A�U��T3��dϞ=K��uZ�������{�ڹ �N���&@�[X��{\��G�a�)���:�77��.�}�~���l���p������e7??7��c��_Z��9qc�W�t�B��T]M8���j'�ݟ�ag?�|�ʲ��Ϻ\^^�@�_*�W��cN|0<�K�?���>|���#��_�_�%����>�� ڟ<��t�lˊAt�d��:�!�Q+q=
��SPR\-�ZnZ���[���tl��|^YPږVg]&�O��K��2��p.��I�,��H�[������X�!��\jt����a5&��hn-x����a6+lƝ���n��T!<�l C6�!��ꉮ�:��7V��J�v׳o��cf+2��pZI#}� �����_����j�-m�V^;M>m�q�e�{u%���"4(����w��N�N��E�(�(?�˙���p	�\Ȑ�3zp,��OenwK��M�tAXWƟ`VW	���u��4��v37�U�e�a�I�n��D�=��b�^vUH	r�!��nGg�M���� S��
�&a�6B�;�I��Jqc+�FT�9Rɲg\9y���ܷ8>�.;�rlA�hAO�٣-/\9�g0g@r~p_�u���I��]�g�2�����&+�(�^� ~H�i�go��Z�Q�}w&����ג�˻/^DJ~���z��'	���=d�ɜ����k័udY�3�}�GB8����`�H}��Pg�P���H��&k\�5j�e��d$\M�?4�e\�_�@i�nq "�h����%9�K�n	I0�aHw�F8��~����m�s_���>;wc[[�E��_��t�������� n�5ϳ��0�b䫸����_�j�.f�^���xk(&@�a��Y$�$VzU�ra1�BI�H��}��r]?"%_Ky �y2��T؀���C]]�[fcs��10TkJ�Tv�1IG��+�z���z��}�D]�E���&�:iӼZ�y|N7�Ƒ�t�Q�B����v,#���|�x��ӏ��O����`�ڼ՟�e@C�����_B�TNQ��r�����:�'�>
Ѝ����=�8���>���&`b���}pb�D���.����k�����fƀ�b�(��e��^��On���F�2S��n�-]�l8�:9r� �P�ۈd�Z!%���{>L�i:V�l�t�������v��JN�%e��<����ٶ�`֊�D��;�(����-wE�>K�i���V-���R�E�<k��R��y���_L(�eH�"�* ��t1��Vu)����X��[�OY{J�T�]��T��"��&�2U[�\��m�b	`������A��e>����m�jšj��ڐ�G�$�#��#B8��<i��8�_�q��1&�~)P�Ԏ��hK%�����U-�~#Z�o[�JN(���lu~���L���vP/�OH�Z͸2�KZ���2zl�஺�c�ڲ3�Z:�l�����}[>�ώ�����S�x,8z��<}ߕ6��Q���c,�H��8l���Ҋ�q�H��|mUw<TO������j�1=�)�Ґu��J��z����=�5=��.~���$r45�D�����4��,:⩂�U��b���+f�r�9SA�ÆF�'��+L�ʭ�x�����ڇUG)P��<�Q�{{
�I����z\�&Y�+li��e��J���\��uA�2iJZ<G1��q~��߄�E�XzH�����=��OY��>:�D>����1��~���p���c���X?`6FdՓ��c���zK�Y�������l��P.b:zD��,��A˸��/E�3��'R��}gg���4~77���",��G�VS�b�
�5�]�ۖ�>N;���/�K���k�\]�x̲M�*h��7 t��X>���}�����Aj�V��@�I�	�'�,4_a������f���ڑ_��;&���%��=�8a�}�Y�\���Zj�/B���:۹N�7J�w����=p/�x����I�\�e؁_�+<y��,��*��y��lKjr�of�T�w�������rO�:)����y:Ci��Q3�uƸ62��7�?M�y�?O�#ׅ̒M������k�~�M����H^�0���I����&:��`<�:N�ܻyl�=o�#~�D�$e+m+M�ɷ�y�`%3R _�/��Iq�:*?�e񌄭�ps�=ŪrӊJ��ʲyG�=Hl��F9핥l��k�J��'=]s��f�{�BU���K#?�A��E�[c����4i�r6Q6^�`"�ϟ��m�h)ƐB%���l��d��Z�X7̳(�c{�\���QZ��S,�^�[��s90���B?��d0T[�e#�]�Z�ֶ�:E?�<�u^�I?~��+�'�����y�L@�Y�����}'�%���	��L9�8��\�b�`��7v�ϵq*��((����sZ��$�S�0��%�oЮ�I)�3x�*/Yvk���i�^C�%�li������L<�U��7L�)R?�����:�	ђ1υ`�1h<��`1��%B��!��Ǿ�[i�VA�����4��7�>����>_z_�L���6&��nG��6oTڦ�	�ճo���Mi6�u6"6x����v����b��8X�t�*���S���B���#,3e��w��i0�s>�B�P4ې��'o�p[s��5����ҧߊ��ˀ��UΌkI4(Ũ}���)7��7��ޤJ���++�j�����A�Ӣ�r)���|�M²�h�1�g�^3a�8!;g�r�:j��@?I�~�f�]V5��_�zր�y�)v�L�$i�|�g���e��=�,�d��cɘ�n��ǹ؜�%Z0RԸ���gq����6�7���4D����<��I�N�R���^��'�~k8�!��A�zh0�DG��\��f#`
�?� A��7�o�0�!������t�֯l�J��l����EYt��$�R�Yyo�w(̨��L�a�ʇ���i"�����\���f��S��)�����7��]$�w[j�`��h�+;��f/'��	�Sr�����p(��Ԯ�e��~��{$3����{��2�v_�?	�zl���VA��U䮹�B�ǅWTl���EqNv#`�2�-Kh�%(�׮n��\�募���U.�x5�_�)W��� 뒌8�Z�57v���`���3I�*��?G���x8d���Zq�T*>P%��#��|���
W8-<����6&ߔ?&�:�
>���Xf�q�s�wUN.���~������.5���H����9�Ꟊ���˚�N؇P=��ٳ�9?&�㩟� ��,�ޣ�Um���#��I]k�hV���lr���G�5|G��ƯE����2�r6@)Q�:c�3&<�k���R�DFS�s׊���/��9ʼ'�i�A�M��p?��+��(1e����	��L!��$�e6���\�3�dJ*;���T����""�@Q�a�i��ѫ�w�.��H�Ǯ�b�$�~".��R��tT���q�J���z�XRL��E|cZ_��C_��:�]��`�$jF��r������>�4:oW�߯Y��G�,�We�#�#I��B��41�[p��Z�H����*�s�7��˄��e���g�m~7÷]�����dG�FT��s8�����rZ�Ũ���c�U�.a��hQ���ᛴqu��!/���5	q��B�������H:l�g��4X����J(+i]87�\xcc�Z�o.���Q�h)�h�����ⶥ>K�!�
��iq��h�E���MgQ��Nȏ��S:��k)��y�yX�].���FÓ���'���RB*n�h���yٍx������u\'^c7g�z�5wj�a����,�7��v��M~��"y�xlr���Ce�%H�_�^?�
I�Td���!�"�(4:0@����x2�y�;�I�T�����&�O�//�Zؖ�F�ɻ1�s0��_J�(���<eAG��������a��, ����3�\�`��2���o�`�v:}��w٣���yq����������գ�3뮘�1a?������3(��Fl��CZď� n8-"����>�t���R坡���J���[���/A�VƟ!�vSJYj��4�;��q�/��_)��R��ϯ��E���/73��_��Ԇ�m�y{ �.�M��	�x1T�E�C �:�E� 5%Z�F��|=�6.����dW?���,wL�!ƫW	�$���V]�mE��mX�F��7��ؿO�'3ߜn�3D}i��!�Cɨ��ҋ"dM䢞��uU�5�뤞����>�٣w!]}����Q��/ԓ����!��jVP/�,���.�S�}G��ʰf̤�}d�	�� ����c�j&>nU�t�佀~�o�63��EF�t��L�k>�-��+~����d�<!V�g�cno	�Y���"Ĕ2c�"H?Nk����Q̵�QykY}s�z�C��C�-�$U��iW֛�����v��5p�=U4��ǀ��q�����qU�q�
`�|z���j,��Mc����h>:>�N|�Y\,��9��=�MW����:�^m�K%lV���X>�����s�OZ7��/��L��G��ѤLDV�+��F܈�2-]���Y�YĖX��,�<a��W��.�:�a8����`Q�_��z�i��m��FH�&��G	��%�Y�>��H>�KmdSPH� FM������V�x���s�˺�ii�9L�&�^"�_�x�����LD.��*����5;�6M�`p<��,�.�V�F��)���8-�,O�����5}]��u{�s���V6ę�cre���Y��@����!�������'bJ��ON�Noc�VWHv�xgD?�<~�'�?�d�qMdб��+F���$��Cл2x1�Hb��ҕ��i����ʺ����;�4�$��p)������������)�6�P&CB�:�[�'�nפ�Ti`5TJM����ą�I�y~~.�ЄCjg��j ��������m�[u�\����]Ԟ?�EU� w.\��s�2�u�J�眃kj�yF�~�L��~��h7�<��BV*���MǺR��-�2" G�'��)fP9���I�|��4��vj� �^���� v��T�~����l��P�~�kZ�����c&��Tr��������C	�媖 ҕ(D�$�fʅ��*t���Zt/,.ZdG+7ksO�]\Tz������*�t�ď�g[Zǀs6;��1h�>#��Ocv����h�K ��`��@
g���&�0
�@j���׶������ �ۻpbT���]��y���d��ǯ/�_/��V�&[?�(ux���]�	EPw��1ųl��h_�U[:�����@n�����BM�'�'�X�Y��3�X�F�ŮDVs�D�.j�]?]a3c���T�����j���0e�@=TC j��`�
u����2˙!v��S�����>�<���z6q��"�iЧ���J�UV؞���e9��e�FE�����M�B�_�%Z=����*e|��Dzy��dU��wY#��73*ɘ@��%��s���T��:j��y�R8pW'"����N��h_�ވ{6'�yeP�Eg����m��z�����]]ҝ�}A�ķ'�׬���ѩܢ��������]�3�{=��Pw�����Pg����^f�g�r�Y���G�����;�Bc:�/s�N��Wz�⍚�Ի� h�yͬ:�N��+"���n�������g��7����W�w$5[P�
��Ã����A�i�C��������E\��􁕨�*F��Pq�W�ΪA�8ҝ�:e�;g�٭جM�^���z��ªcr/{u8�ۛh����puq1ek∵
]Dl���:~*ZO����z�YF}�:�a>���]2p8��I��qحp+��0ְ�_�/�V��x���}�S_jX��{0C��ԅC&=J�$��Y�)��K\u�f�������\+����B2�ese!�_��)�dok�F�?ҽ"03"	Ob����m�o=�#��v;�˦�J3�TE5���w���L�V���4�,_��s3Z�\�d!6�0���Y�#+�O�����8�Ɛ�9}��3�����Q��qU��R��~*�$r���`�5�چf�Sִ�e�G�Z��F������P s(�}V)�흪bׯ-�[n;�yT�g57��#��{����eu�Q�P��c^��ϫP��X���CZ*�s��������~U��~�8�������7Di��ԇ~�Y�ض�Ra�>�������vL�o��������-H�����_+��{
=H�����.������O�{��H�b�ya�]�z����&�UE\r����4��1஋��u��*�h���w�r�BV�&�PʚY���&�A뛛�w`0��P����5 �DU �#���Y�T�KՅ��#N}?�۟�锁���������:�������� RtE�꟠������*>j�ˍ�Sy]!L�>������-G���f�R�=�B�QfBd����:z���?M���'��i}[$tP(���|���+���j9-�e&k��צ/�A���--���P�Ozӱ}���cRd$
h��4�ݡ�֕��63�̣���*�;�/��� ����@�*�o?%V)�6�Ľ��믉�u�H}�q㇁�c7�8�Y�݃��S�X%���0f����v�z��Ű��a��⾡��G�P�%����_?�T�n�I�R��v��CѼ���o͚	�x"&>����T͇�����+;|^\���3���ik`K���Uޕ\���X����+��it��\=�� 
/��7�!�"�1�oї���x�'���J�2���Է�ϵ���uמ=N9jܑ�(�淆����\`G��{���ѓ�N�����9@{���N��F_��z��ƹ���s�Q㣆�ߑ�O��Y=�:7��������n�����݂�&�u���r����s+I&�(:�h'O&P���scN���1��{_cj3��ُ��f�"�fh�)Wؤ�i>�X ��U��������Y�_!j��po����0b�m5��-�;u\J�.���G9A*U�w���݁�ԃ'&��+��أ��ҽR�m�v��=QS�\`����ԦH)u�UƮ���d�wa�;l�����\��/|�N��s&��D�c�G�����̨�z5�Wy�kv��h`u�υ��u�~ڡ�86��2����b},ނ9���%��x�M�r/݋�(�G�����x}$�n��hVc�#����6@�d
���d��	�N�k.�|.�;i��+=X�V�$H��h�8�R����_����I\��E��y�K�M�3��A�yʺ%n��q�q�I�:�$/C[��{-�T[|���P:�ق���FN���z}��������ۣ����٘�,F���N�X5@�X,�7����B�-����-���ǻ�K��:�
������A4B��+���@��er]����V�*�:��X9;�鉈�#-H ����e�>���š�<)��� ku:��/���Ů3K��~��V���'�R�R�:<�VW�J%�jד9�#r��G�bd��F�7�R�Ï��m<�\��P��5ݸ��'�4���y7]�8�r; ��9}'�b�+ojb�'ۆ-��8ӧ'�HX�����p���w���{�̔�H��G�ܐNG�x�yd��D�jլ�����d� �Y�u��/&�~��f�{�^�=�/�I����ԡ��O$M�2��6��_G��ʵ����""����@Y�d�v|� �+��U�'����| :٘5�
��s��Q��na��$:'r6$^L�57ߌ�|_�ڋg�4�倂M�I�6�w#WC��]��$�{\x�l&
�.�<���o>K.�|}O������C-�����o�`���5�<)�鐹�(�d���\�\�6�w�§|Y���J@���ܔ�����=BF& MFO���y�����(��R��.��
tL�A;�[:�r}���!�v��:ţ�&1uT�3]��	�
s1�/�.���[�L�5󤯺�OE!;._7��n�5�� ��̅Wœ�0���t퇿LfKSם2�O�(�ieL䠩�s���t�lY�!�x���٫�������~oRP ;k
�W ���#UA�\�[�@���帺{ˀp��r�"�K5c4	}_e�������7|X2^�a�ZT��)I8�ׅ����-ԓ�;˘L��T���&*Y'o+O��ͭk,���9q|j�zi���f�����;q��1w~fs����~����ᰵӵ�bң���o��(�^�.�! �J� ����UJ.#��m��YC��N6�ј���������:�cz4����-Z��Rc��&�����<�/�?,,��:�w�F�~��mh�s�?q��tq�|_��v��dխ�}����z����X�蒽���)�)�[�-pZ�󺚍,�����)~��!Y.��gCe��Xv�Vaa�&&F<��qqq���s\�rl���x�2z���'A����A@y���ǵ��.��m�-���M�&�B�p��x1��i�m#�{!&W@����}?��//Y�ju��i�U=-H����kCoں��1������j=���[�g����IO�&�8���o�}��}�/9~��8D�����UΛ�J �t|���([�*g֏j�l{�X�jP���7al�3�U�u��u)K89k��/���)��V-��r^b�����{���S�c�6|¦�Y`��M��f�AF�/���ET���	���h����g�U��&��_C�Db���y��!ł������+�ܯ����͚t�p�#�sP��=:-�[� e��0��fV��W��Ll��':��S-C�����MR�;�����yN��%"&�>�%
�� ���I��}����!$V��5���;<��$�J��nD�|B	Ŗ��2��J�x_�j�:�{|���{��%��jjq}	��<H3��|[>n��/�sj���[+sj���j���L%UD�J>�\_+P�! s�Z�撕A2P����~~����pL	|�s���f���H�rq�9�����GA>������T��� �[�ޡh�j�ݔ�Ԡ�|� �4�faAͲ6n0"�e���s|��D��k�x����{��� bj���ۋ�?l?wH���Ag 0Q6��h�Ap5EMb��3�#Ag&w�����qB�m+TB�,Zu7\_ؿ�|B���W#��%q�;��|/�b�'s�ț|�}�x�;[������G�g��o��d�V�|�����=�+1�ĭ��>�<�8
�"�9R����sr�
�u�"٬2�];ߏ7[]Z��y����6ߚ��,|���%���E0;�x���/�%�-ͅ�x�&�����v0���蘭�������a��;6S���U�" �3���ЗҷѭΖZ(�{�P�G��rá��y/J��K�:'/wO�po?Lf�Á��{���ߖ�%e���!J�|k'���:��H�'�c��l맇��<f3̔�wk��l���x���ʜ�T�1C�F,M��ؠ6v�2�� �� ���*[�OV�%�~��qts��Aܞr�E�t�u� 5�����=����뇛�To��ݽ��%jU<1S�q�;��A�&�;g�����l�7�RB!m�ۻú����]��f��c�=� �A�F��8F㑝�	בee��1�"��+0��0"���Nl��C�׸���������g<��wt��Z`���\C6�f�E�qRLf�*��.����y�_z�W���<[1�ʊy�n�+Z뫔\���.������һ)�F�O'��G��"�;��Vᚓ�z�D>?���)���Ʊ�j�bW����;?��B���T�P_����_�r����~lL�x�>9���G��b|���J<�G �}�~���0"�H�C�:��ƈ�t���	&�Zݼ����7����H�T�*==ͼ�d҉����[��P��G�<_$#A�Kpn��o�H{?-6�P�x��-zN:��Z��xtO(��n�$�d��<�,�̥��O���gc'����O�z4 V�ؓ� ���9�y��~��3�����[�n�h~��Н�0m��]a#y�'���sG�*۩�xH�<���5yy�磍ۺ�qh���k�Mw�y�r�G'H�d�lIѫ���W��+��O/��j���P�t>[|j'�ҳ�!�.B=�R#���Hâ��_�����g�]�\ܕ��'�٦��K2M�-4zݕYy��}]_����H�q�C@��~��ԫ���s�R^���~ϥ2�ԩIOe&2�h��g��B��v�G	�М�S0k����[�اo�_����-�2����ˊ�WW���f�}q@������	�q���J�A��n ��(��6V�����}҃2�}c#�'�ʖN�5bݵ�[�ٯ?�{"�� ��"���1��������VE��> O��J�n��
(
Sg?��b�����푫�'abb������1�r��w������`�������V��D��e̛�����OmP>��I�Ѯ�E1�i̓nֈ	Rk��h�/Tâ!�����em�¶�q�G�0�>Y��n1�U��0�X젝���Lnm%F���U����}Z�)��ɀD�ݍJ>υ� zM>ޘ��Xq��e����m�ki��w�3,�}�����t�u{(l���U���Q%�u��n��bd^��]t~!#�r(��n�~����T�Ul�տ���xZ�M=w#�{+�r�s�c{9z�}/Ûk�����8aU�0ĝ[�L�S�Z\c�3��	�ޓ�&��7n|�`�������u&���a��{ن�J����JYek��3~���f��΀FQP^[�l���������jGa}4c9�dϓ5��ۮ5�f6�f`����w�2��I�؛_F;Nm��@�����
�*|��r��U��M�D�|ԷdD�Y�WTR��"яS��XJ��̎�e�O�D�_�2�(�T�J�1�|b�J�z`"��������\�me�WhD�(F��b��I`�Ɇ�f���	������B�Q�Yo�=Q>,�Yܹ���=��;�r]��^�.AJb�}H��O=�������n7��i��m�u��o?ڀ��U�z��';��S��o��@�����o>�� �x����+@�7^��5�]����qW��4	��dT��F��;�m��F�P�_����^��ݎ�K��V:��#&x���b�>,��Y���&�� J�D�ލ�x���p7a���X�\���+W>��T-R`��O�y��G���3-�4�?X�X�DKy���J�Ϸ�"0�(�uv3��e��")P�m���:q7�͚��Sw'�w�ƭS��hFO�V!'�M�5��S�ޕKZ?�3|4�ղ_���M�]��.0x-^__{_O��WI^�K��C��؋��cxU]��a��wT�j�E���Y�M�������Q���		[Y�E?��>e��H�L��nݮ)�&Λu�<����?�Zt���ɨ't�ᫀ���}+j��4e�G$e�A�#��=���c�_�p[EK�YS�0�Ms�k�W�b�>9�86uXi�p�d+D,�J�.��_#�%q�S�W*0PC������t�m�ڛ���m�n�����"���Y�J�%�zRN`}_J�>0[0A��!���h�ݮ_�k5�J�czNڝO>g��G]��@�6��e,	��g'e�*\'�b�K�	����j�!�Y��җ��d���޴{�
+�x�Mnx��s+2�	�G.Rtb�������
[�걊�W^C��v��-��'mwA�S:&Uh8�B�]��e,*%�3����e���݉�Q:_�!��q>wc� )��\�:��dok�YW�;z��5����#�> ��_���2W��"��l�2yF#௎����8�(o��ڻ�H�������=�wdڎ3p�w�^gn���'maK}�Sg.����6��'��� ʴ����68�v�������M[ ���	��í�DG��;��Tu���߸���O���0���%6V�3�T �[Bd)���o��7�<�P��{�1�X�R T�ov��zXt�/%n{b�
���8{Ĵ����A�֍*M\QǛV8�6�Q�B�=��l1��|���؀V�_�m�e�++UpG��g��:�������n�=�@U�R۴y�GC����~[ej�U�p�(��~ ��v��R'go1��R�|B3`������7!��f}܌�bv��)WY:v;�q�k`���T������^̻�5�uX���E9|r��� 
���Ҍ�-�N�e���T�n�c��­�D|�.��\^zi�![���}x��eVj��!�Y��G$��	V�?~��,��j}�����́t�������9^R�����*�ү��!rN�.ꟼ,[�ɰ$Z7^[���~�/R��m�����E�q�ik{cw]�v����,H@����V�����߇�L���u�`���۔?�/SS�`+�U��qr�r�@˚��b۾Ի����&g��o�4�R��e(sX*���t|��ͩ�y��/�N֫�>�>H��=��zouؠ��!�U����=�J]�(�#�����5��\؆l	Zj zu �����z@��8-�����_ڑ`�?OE�x���S���M�G*8�_X4�=���{��_�uj���D�{�=z�\�-²�l�ҫ�N������c ��������4�{�*.>��o�.mjnaШ򜤠�|���Ɲq$���h��iikK�A����gރ���
���UI���TR^b+��F�@W��l#x�-��)wu��{6�j_ܑ��m7��r�J.Nz���T�Ҩ�F�����Ĥ����O�?t��Sp�h�Q��~�BF�?P;U� ��բ�nF:ݶܳ�ῦ#��L+@u��8{w����������<���-�N������̠���U�,��PCv<d�g6������(2���:�,}"��A���sG�����~s��v����FHcީ��uyRS��ia�����V=L%��̉�#fB'�`CCJ���|�Z��mYl��Ғ����Vc�!��������H��o�3h�"���?R!��:��X���g�D߉Xճm�`x�/q*��^�t��vM�?T_l�����Ը�-����"̖���59C?�D-������Rt���x:Z���5VC	����Kx�Y��/��Ǚ&N]��r3{�Aݨ+�$����:o����ҠM����CC��]$A�'�ǆ�f��B6L��li�� &w���54u���������a���̓�Վ�2�H�@��~��g�]� �r{��T�l�%��� �����l��/[E��ث��	����<UBda�=`��^eY3�O�6������V�^�]��s�"��XN�^[4����&��V��Q��B�\�z��g��7� U�\��	{࡭�W>I^�KW�pR_w���}�����Æp]��˜�"�o���6A���V��i6%r��u��j�I���{H���jWt��E:��j�--�|�v%D_�\��z�A:�d͉!w�����{���~������U�=g�j�
�*ꦶ�NGE�/�#�ۜX �'L���IN�s��/U��d��z�K�{��5R����4[�y������ب��&<��(4c[������,/?�x~�5��;�+��N�]�bѯ_{�V4��T䵇��5ʴr���T;fB�TX��iz�Bߴ
��y�*�,�hľ�κJ2�
YL��>ݠ��瘶^����2��=��o�q[���'{/�Ai�������N솾q�_]�& �_���ڤ�c�U��hvsޝ_\\MUŭo�8%�h��o����_eeH���.Z]e;�g�p|�a��� ��� ����\M!_�������W�!K�����aJD��j�����~`�[��<jyv�^�&���7��.F�-5C����n2�]��FK�$H�^?���@�\�� T�{�4O���S�|��7�9��:.茻�?d�N�0ڄ@��>��QH>\[M���>�G��O F`���cW�ݣ_]Ν+(� O_>�&K��'tqLĮB���~R�L�#�2z��O6��\ ]��>G] �$�gk��1oj�wה�q)c�xh0Kǘ��%��<D�2UPZ_h�?�zIHF}�ގ#�fcc�����a��J#%������<��	Hg>/��"x
�wA�e�T�쭑z�r�i6Ѷ��P�]8�b}��
k,��j|��#����%Y�o��v�''I��m���3��$���Ř��}�3vvs)8�\�'�xֺ���-@��e-Fih޶�y�����=��O��� {ʓ������.g��g�(D4E^:��f���z
�����mv�������[.�	�A��w��q��{�ڧ->!^iHw�Wc�p��.���$^�-آ�����Z��_�|	5���Six�偖R��L9����a ��m����y�!Z��ʈu��,�짂F���ɣڟD�ò.s�l�4|�KU�|:)��*���~�!TI�E8	g	S࿐�;�t%�ҳy}?��{�A�����?:�|[����	o���f?t�s�"��$�,|�[�I�kɟR(6o!��F�D��[[�����2�8w�r���[�16ֿ�ԝr��k��2�ۛ��8吗��~A�{{�]ˑ]���7_�@6b���2�=F �O��D
mi�bL�h�E�n�������K��A2�ź�Q�7*a���dE]3f��&�%����y2ݤU���X��r����oG���#�N%#54|�S�r-�|tLQiܺv�����t`fBT�?g�<e�����֎��^�*�.݂��ӻ������
���u��Nh|o��8���w�9kĺz��q��Scՠ
u�m��X�����$���Ǡ$�4v�L�S���p��(Dhlɝ.�����X\KUZH��i�	��P~7�)���M�$X���|�~PY���8�J��wA��Ҥ�0�F:�n �y��=��)55��rv²
]y�9L��
U�l���g��1"�u+u�_rX0s5�c6��m��ݯʻ� 
�%%%��&�/�SQ�C��l[��~�n2�{�-I��mj�I�̕*�0kD���ѱxn�*k^�9�Y��>�B��	_�`NX�;��O�W�5�< -���ty�3���t9tCb`���2��^�^$n�ؘ��6���� >V+����d6k��C���[(�q��&%v�Nb7���z��&�;'V��~K�DULH��7,���oޤ�6��朗��>���gm
�J�R8;��R+4�*b��8;�cXb�EGG�G��;��^��|"�����m�o�TU�Ջ�"xzA��� ����|� ���O�6��n_��v��i��2G���s�N����Mj�,�\��`Hʥ���l2�ܜQӗ0[�������B�WV���w���������pw�<��Z���^�M�r+}=�V��c�.lgVf2��Ƿ�*v�o�Ѕt�b[��+w~SŇ�8��) ��Z�C�g+������f͛L[f�G�P�}R������<��뛇�;Y��WC&�/=+dN�-].tWĺ��8��'��$^�Vˏۮ�+-���k��?^2��)Yo:zq��uN{tdi�8��+��xf�$T��I?���w,y��������Vű�^�ԙ���'���i�Z<����X�g!ۄ�C�V8F}�{�:b��Y��j�#��d11��+"!��FxW\�e-~�sX�ǩW�(�xss3i�3;+���6w�&6�n�M�÷����iҼ������^IvT90��m�4s���G���zR����x��V8�PgX�������:��J-���rrrbj��o�׺nO+핛�/Y�<2zL�$qZ0�4�#�>�⇗��R	��>��K�4^^��	b��
�Ig`7�,�r^P���4"����� ��z@�A��lR9��/%2f�v-+�u�on����U/�{��%8�����]^Rd/83I�J���.䊟�
dr��I�w��
���I`PBU�Iۡ��9�a�e��[c)�/�a��K�Ipwo/Ɋ&7���#ר�HL ��r:9w	�ޚ�����}�d���T���Hg�,���K�ϕ�&��W�8��L�:tt�d+~�S48�6	�9��[&=u�Tk���:�ݹ}�H��h.��.Ė�]�S9���3|�8�
RIfP��̝8>�����ɺ�u%�j°�63�l�w�*������hp���[#���_N�h��t�8xR��������o�����xW�K�m���Z��H��� '��ѿ'FBy0�*K�A�&�&�W��]ʷ� �U`߄J��}1����xŐ��*I��M����{�Y�T/i����yC$�jc؊�F-5�ݿ�kE��:��T�&n��������ɢ-ƕ
ɡ���W.A����z��9�Y¶�/��T90�g�����(ظ}����X�~��a���~G+=N��)[� %�Ł�/�����7��\D.b�))dp8<��ar��x��G�������'���N%u��ŝ����v��cדt����|�.�?�Yć-s���� �!���\����g���Q}��7�|~����W���x��{��ֶѳǠ��F���r92�����,E(r]r�<={��%0�PQ1*��=��y���x�(��4����j�ﲵ��6�m���0��b�ܭf��-`D�󁺋��l�"g���Oi�7�%���{vβ/���P�����S��Kw�������1=�06������)[�����e���1�*���;�H����IƟ,���AQ����NWMZZ��$(!T��f�1�}�?:;K���i#��:�"�hlT�'��z��p��s#��Gaím�+�����YU�����B�:�H��{Wս��.;G N������	z��qt�aQtm��I�Z�%�������;�i\`��k)%�Db�%�%W@J�}��g����������LM��|~S�-{��F���sw��$�Ժs�ع�bi;y[
��^f��HT٥8����X�a<C$�����u\.����{9�	l���p�����UBI/��|�i�aj��jN�7�������x�\ν���F)��d*$�e2�M� ǖ�A�r���EZl��o咡�eT���
c�"u�ϵu�13�Y,�l�Ґq�H��t�߾Â�]�����ϻtQo�؋�
�mEn_�G��m���Cye�*� \¿��М~�:��V��g��&+�L�sIg�����9Օ#<%���t��4���Oǃ�~�?Pi�}H�Lu�oG���-������֮�!;�{���S�Tl����$D_ȓ|+��а�;�X����PM�p]r�Nϳ���w����~�\��K��;݅�bq���>���&֑���?��&���%�q�6".2M;�׎oz�P��h��g��N�FH1�Z�l�m;�VJץ�� ����W�J�%F%���?P�J#�tC�����W%o����o�@g*t��/�((�UȘ�j��?�n
��XL9|������␣\���b�������`�?`���ɬѲM���>�)����B�&��n/�<:ڱ���8;�ů�	�g��''XO�MDmrHl��<

[���lF%A��+�~��	�okk�/2X�$���D�BQ����={��;�	j��M��L'��qcG[Vr4n���%p�1�Uodqս�1�a1�}�:ܴ����$�l&���i�˻E+O�s׿���x(�e�|��0K�h�� #�Mv�c�9���d��G��+�ӯ�'�~���\觠��:Һ0Eu����`C�Q���.��G���J���8Q�S��7eґ�e� J<��ws^^^ݰ���CQxx8���b�\1��@�:X����s�U�����]�.(jp�Ĥ)u>!jpe�Qٌ��9�6�" �j��@D6ш���?����gegs��n��enK����Ȱ���l�������P"G/��Z��*p�ަ��ٔ�����>��ʪՔ�'�f��e���E��1u���{� �4�p:��f�x��K�uӿ�5�IuǴ7��]���ҿ­��K\�g����0�o�N(��b��3O��_�8ϔU��Dߍ��ٙ��E����D3�gq�k���鮃��M�^�H,�����WԒ��xw�=�,�^ 02��e�m�w���gzOҩ��b�Iv�]������7�{{���KN�cH#u6;���mݜ0���߳��9R?<D�0���d4!x�z�D�(�ڋ�@�B٨�DDpp��}��o۲����������� ������W������7N�����89'�Q��7�w��Ɠ�L�����qb�f$����fY�{c`t6�L:�}�$�[B�>w���l�<��1j~�m#PQ��YM,m��*;�%�JD?9�^D�ty{��K�F<
{[�@R�7K��s������z�<)�(�r.�*>�8�Ch%��>�u�j�U�J���(l�:�yZ����KJ.q�K�ə�#F�]hf/��p�填4v�ijU�{ɳs�1��xR�,���/�q�B��~n��7����uP�;�PZ�W�jEX�Z�/����Ά"`��+�g�|p����l�<���l��)��]P���ȩ�E��-�G��ѕɺ�}��N\|K�]L��]=�Z=k)�M4<�a%��7껫}�$�����pw���a����
�\Q..�Կ�2%��8xg�_Ca|l��č�Ǎ{�K쁛Q~5x>�nl�$PjC�J�@�+������:7;2O�?�µcE�/��$��X�:=~�u�+��0��4�55�k�tn���H��CXGk��t��ۡҩ��V��#-��y�Nm�>�,$Y����W8�ax�?-�����GG����G;$*���d3H��������*���Fwܳ��c�e�gG�<ۦb?���V��6;���w��8��ꁰy�����"/>D]A�
�#����(7C m�tɻnJ�F�M�f��!aD�D��0���e��
��7@!��,7 ͉���s�.��'j�Q��*	�=TP�,�P�~��V����@ �tzǀ��{֙�/$�7 ���U��)q;��%���"fo�eC��猋�{ GP��nz���*��q;\)����Cx 1�v�Z*��Q�U�qj�F��QK�U/k�1_ߝ�N�F�z�7*�,��b9���m�TJ���d{��E���3>^7q(�;�sh[&��9��M����G��2���~M�z�]Wy�ߞ���j.ӑj��4�=���	�F|��DќM@G��i?�f���Z/��PJr��������A̩(`D�����LT�݀�yz��-�+	jo~�a�E>��j�s�Iu�o���SmiF�f)0��O�`mD=L1ڬeC��A��?1�*��Ra������2i�Jк�K����أ�Ԩ>a��d��:rc(>��48��O�n�Q�6�TnqRqҙ�HP�Uz�h�gZ��X�o�_w�2�۔
~�vBFEQ��s�Lj�7s���f��/|IsXI����^�c�F�ri�q��'��}���I#�F�Q�K�i������1T�X(���x�MN~Ng���(D�W�?��/��G�v�{�:3^\HIoo�K��ONΤ�E��5��t�?ng��xS��bۅ�23�/���S�Fj@�X�'Ői�-��9����<��n+�.��Z��l�.���5���N�q/Tq������7��x�����'���H�����W�Zf�W�&cdA[YQM:z���(l8�����0�1��S��a������Y�nX1�I+R*]\��?K��t�+S^P��Q믓;ʷ�Q�ݿw4c�KV���q+f_ P��������/��/�v&�C x��f�MZh6iU���S�E�*7r��I���ҡ�)4"��2�لa	K����`�D�xV<U�q���1Cu�u�z�p�������X���`�KBw#����/|��&���@����i�$������x+YJ����5���f�p8���=�>�a�2��:i��Z�3�[ǝ��7�mLt�l���|z��g��:��1ה��r�O0l�@��d�&�������H�e^/+U2icxQ([��JǪ�3u��`�~�B��0����,��C�w�[�c��@RzY���˃�3���"n����m}�����!V|�0����U��M�[(�����%� P^<��V�Bc%-���e!d�_��;dblF�9�9�lJf��q8@����SD���E�<�I��2�R*�6����}c����˽���S�*զN@%N4��R~��k�t���)c ��ڊ�wo;�����Q��4	a޹��q�Y����A�����0j���_�UI~YQ�����u�}��a�T�cY���7�m3ϖ�GX����7�G7l�j��'��-ɰ�+)�&�`;����d�Pv�9ˎR�QE���2�S+s������.Yy`����}��f�חя�����\n���5�_�p�8(�
�ߞn�ԫ��2~K'�E�鉳�ʋ�m����yY��*c*7e:�It�t�aa�&o0,I]�-���I�Sh���@J��]n��Q�2����)�z�	�K���������s_�������l0(@uaϥ�e�i�P��h�[��v��̸XG��R�����K�oY|�v1%t��Vm2�	7��	�D-��i)�Eb�y�-���*�D��m5�zL� �d���GM�b������շ!F�K,8�ڭ��B2�-�C�U�)���^�&PmD"r&�7��%U۷<������2K�IΜEX��L[g��w�b��	�ظ���33>�%9./uΞ䲲����P0�9[�ttsc
�0*�t�21���+����5�j~m.�c+�$)v�v.��P�_�M��؇�k\��|䢈v'r���:�������WP]�T�[tc�Y���.,G,P���Ku�����v�[P�p����ؿ���7��Ѷ������q�S�)���9����e/Ϊ�mn�)�f+�VQ�O�&�+˶��������Ęȳm�����.�)�dΦ�MZ0�m�,O������%�cV�zP+ ~��3����i�ĀM����7fwz^��]�N�������%�,��6&�vy���µ8�Upˋ�Mc���0��Pl� #=*�	���hgg��O�#Ğ�x�$m�=�GfR�	.CQ;F�H�U�`���N��M��"ZeH�6�(himy�����P}[[O�t�����&�F��]�*�y�}��%�hi��p�)��an�a�L�29[��z�Gж��u/??����=+~|����<AoiB7�}��B�4qu%܅}�G��P`/�"����xn�m���"9#.%�D���ֿ�2�`QT�U՟	I���G��y�]��a>�\_�t?wu9ĩF݅��ho⌍�H�GW�؊___cF�v���t&�,�+W��o1J9u�Ν��ΎE�(!�
>(��%�ذvӜ��pV�E.��XC�Q�Z���F����G���J���UCԦ���/]��^���V4?5Pk����ur�o�I�ߩ�(��J�T]�H�����J�E��D�x���/ԕr^�e�v7!N�zנw3Ս�C��Z�U��).�%�.z�.w�d�_x�jd��p5a�����a�f��u����v�iҤ��-��}�U5�f����P��~y�e&�Q�]-��G����!W`��J��>�TE��w��O..�itk�q��u�d�\aF�@a#��P�eZ�R7��c��q�/��|I���Jdl��kk�4�d^P�U3�>*�صl�4~%}q1��`�:����'� {��#sV}��#k+ͨ�g[D98��2�{���qIW��St +r��o�mY G	�**c�U0(�d+ӟp J���q]��)3u:�G|[��NH���jw>T�MO}�����l�]�3���9W��#v��j�~A���$���4���R�F�����ܿަ�\�"n=�����K�{���cX5�X�5S��nA�v�ןH�H������^j}= �Yj�d��,pkb?J��Vh��wL"��O���A}��>b�����S��s�=W��F��ny�	�%$����{��*�v� �g�-�l����#D~�͒`ר +*�O-�eV��!�;M�T�2 Zˍ]V;*2����@�hz��ӥ�)M�D�ڒG�%u���v��ȇ�c�R�bN��A�`��)����Q���Z%^��}muJCs����-�C��)�l#ꂠ�3oD9]|0Եswg>=���Nz���TM�������������e�Lۈ² 081�z��������W��U6Tl��I�a��4�r�Jƍq��lBp�}2������X��{���n_�f����;DǾ#(ה�[��҂�~`w�6k���_��i���)�������"*q=r����V�Z��,
5��е��iY��|����<��:�núQ�a�?�����	��@y"v�k�܀�K�������Ȯ���Z纺��#����^�9��Cm���@�\\�����1��>��B,��W9�r����-���Q#�q�P ���Jv�W۹d�g�,���k@�0�VI�i���9K)�������*��5��Uc�)@�5���]oV �0��q0����~%2�&Ϩc2�Ɨ|z�&�:�(b����i���Qm耨S^`�2'JN-�o����J:t��/@X*�i�͚WO�)h�D蓭���`&~ܗLK"42]8�T��1�y?/��̆zL��L����� �	�B�������7�U����I~SP�%�'�9��)��i7����ro1m�j�Mv�6œ�ٮ��2�f=>Ez��;�qG�1���zO[h�X���Є�"�ұ������ޠ���y����^�в9䭃�w;qg�҉��i�m��u��y{���ڝ5�GXd�U�hc��|Q���)q=��U�����O���ʟ.k�&���Sg*3_9*� ��߁z�I4� J��K�[����32w;�췌��$�A���Q�h�퍦FgK��
�%
;� jAjdP�n��ٵ���d�
O��YX�fi��1���^Q�˶"�#������МK���5h%$$�Ѩ$��3v�dz�����2��QL���/C���׭ �u!��k�n�1i��A¼/�����㠯�Tw�}Hjø���ۼ���������.�֘�@H���	p,�EH��ad�Ǝ���8r���ݱ:�3�ŀI.��T8�o��=�9���{��S����������ź���tU�Y�,ׂW �xS]��ݟ�:�x����i}܋�ܖ'����M�KY�Db���1� N=�A�M���I��G�S`l��˻{��ܑW�L���s;�yk�!�*�Agj9�1e'�e�_R"!�^��"Ũ*���DH���-����]����_�6�5�}�F�U�hD�-���@Ky�I0�:)7p���P'�c�i8vfک ^�"���z	�� �o���;y{�*Á@x��b-��.���r�\�tp]Ob[Fq�Ճm���KV�V�:E��
�D��F�8��SELS����i}�u�5;�̋�ӨЛ�ԫ��/ �>���j}7\��4
��-sti_ -���[�]۲@����J�K�wu��h)5��ʚä����**�''?���'*���R��	iY�Lя1�ka��eI+4h#�4=���q!0���\��;���TW�d�E�[Ɋ?�1S���7�z����;;���l]�Ƭ���q�󗀋�M5r��0o"�b�w��yeLG��	Z
pYR������݀4�?9����N��S�ߵ�%W��:�[��[�͢%�2�;{wIg!���c����=ټ��[B_
���̼|�������_���-�[����<�^��*�Ĥ-�F�6�ȵ�:���R4!Э�;��n���L�~��c4Q����]���?������i/;�	$З:�pހ4���������Ĉ��Ӫm9>ii��	��z!Y��x4���(<y���D ��s5���k�2w�uo�}��� 
���!Ʊ6�+=�Ҫ%S�q���Ϲ��%vٔ �Pei���74�
���r	dq�L��З@�_�M�_���	�O`h�pf&��*���!e�%���Y��XC�V�79��	��T��f�B���y�W�ZZ&Q�6}��kQ�m�:M*p��.E�7$/
!�r���D����%_�������S�+q�7�4���o[ݼbA�6e|���u��s��9�2��.�GNB��l�qD^�h��K���gm�R>�\Ұm���P���;ǜ���/���O��#�Xu$gش�Y!���m��E�\F�fAg� ��"ED�B
�����ub���L��Dp|P7G3�#�PfA�+��kV5(�	a/QJ���Y� ?�o�S�ds���}�ccc�����[��������0��iʙ`A2�xK���v:S�k�	�Ԁ�)/mZ���VT��>�����3�nt?������dR/�j�.4���Ԙ��"�4.0��#�<L�:z��-@�l����А4��;��������*.��C����Cop?�6�����@
ޕ����g:|HKC#���E
�v�(V���\��F��(�z?�C��8z�qU�z��u����a�=��}��n}�}��M���q��'�*+�!����s����Ce�W��K\Z�K��[�0| 9�*�Gә������"Q�� y~��O��n���/��-�/�?*P�T��:7�WI'q,��+�}sSt��『����O���a7��/��� ���|M`}�+,T!�	�
\_�Ǔ�n96O������[���W��/�rbU�����x��:�Z������A&J1�+Vi�:�����!I&m������g�����N%�M1�Gd�J��6��/n�%8M��)|g�r�KV�(��B4٪���o���!6d�N�A�����n�X�%Y��Ų�,1�*�w�@�s�'�,$\��}1��hPg&Q'}�����7U��R�j���h>���Y��_QӡH�)F�垷��h$T�U����U)��J|��+#ʊj���P�o�={v.���@�\��ȏ�o�ۑj��1�z��^JE�s��\ Y���X�5�!I|�1��.�,��->��W�o>����"��[}�<Y��^<Ht�҂�>�9Ol�5�$ݕ�E������x�%d�U�^��|�c�~=Zh���tZծG�Z`�?2X	U��ɚ�5%�C��~�^]����A�V�Di�k�l.~��ʜ���P�C_�[�x���x���G{%��J���@I�	�؍���Dӂ��C_`�"S1;�6�����J�>?i�/E�i^)��hЙx����V����R�l������#T-��e�@����C�0��0yt*�T�00�4L_k_ܑϲx¡�ӣ�B.0,��bX���-ޖq�c�e<=��ۥ����X�}��3.�.��T��ō`˫?/��󍒐⿌�r��R�b#VQ�_:}5~^5j��\azn�u��o���:��PjPe+�&��C��p3~��쇯bP^����Q?�b�%�B�Zm��+�Q0��.�
G���I���]!`Z5��+jb�Ȁa�����eR�_�l�w�l��>	ϔ�쯕�F<^�<ܥ[���k��	����1�!��su��c�g�jPJ5�L`HH��e�W����,�55��I�)&Z�h��� ��������*T�vP�N9g��5>�rm�Z�m�\3�n
������!D����E�i�޽�����a^�I��*G����&&�@���_ߎH�u�+4�2F?�<ݹ������/OLjܩ�f ��Ћ�8�kQ��&ؾ��[�>�E����"T6_��{���"N�$�8q�I��Y:K2I�R[��k<��x� 5r��AV�\�ۃ��U��<{�`�N���'���I����E�]j%=D��	���]<��-F'ۧC�'ݡ_.j��p�W[{uヰ��w�;H�7�(��/{/ee"S��<�V;��1n��h�Ji�����*��������Ÿ@�߂�Z��>{ ��/�+��~�~FUJrrO]:=-"д�8���;]�Q=�Q�㶓s6�� c��ӛø|��ORZ�@���>�6@��w ��`�i֬Q��ȣ���2�&�3��*���BZ�iME܍`�+6?.DBV�u�Ԋ��uԎu�ߛ���0Zhp4�Qܺ�ϭ	FkQ3��*L�yp�x������s�����Jvs�2��l�d�$�)��s��G�7��~+"���t�ok<W�z�=�b��Dɖ5��|�|���5��Ť%����"+�d'W��L%��J� u��%��	���;��nک�ˮh�ʏ��5b�������+�R,R̲��tN�,q�g!o�Si�``�s��
dS#E����Q����]�އ�b�T���#����G8�kN	x��`� �n�>�׼�`���_{��8� ��끄�����h�X�#G������}շ������q��"��32%8\�2O��^���_G���/ԭ�8E-����'����G4�r魋��m�r�>~a���m�S���j(ؑ���R)�&���=�6������.�#�u�*���mFz���d���+���G��;]��4�SAj��߆9GZ<�wZpig�%$���L:3]�東�q�a[�k?$Њ��l��Y��g�RQ=4D?��;9����BSߍ���Ȳ��Z�[&?g6ĉX�( �F%z�|P;�ekix������K�S0ב���q�6���n��mbt��	_Ҩ2W�#0�������+H�����饤�����.Jνp`���ʹ��6��3�_�)W~��=`�ߩM�%PXf]�U��X�X���C9�����K��`(��AF-��{�����FX3�ޝ��	�Z�CT�n�ĕ$Ѫ������k[LY�'�E�j@�}�.������j����N��a�`ϲL1�DL��Y�e�;������v�=4�s�Fg����C�|^����o[�#����k؋�l���ښ����;����}3�Η������U�:idM�b#ō�aU�(<XI�ZQlL	�~<���)hTI�J�����dg���D�|��.����qx���2���;f(�K��-\����j�yס�ҏ�ncJ�<�VN�m�C��X����t��먲^�i�C����XL����SX�W�~��|�cTcP�30�0b�!eU/m��W����kC���H�X�./��I�/�smMx�U��h�ŗ+V�����'0B5��礫�X�M��Z�j�'g��3H�T!qL�`�Z��̀hJ��ϟ�-�* 0#I��ʍ;��<)�5��9h���Ŝ��ӆ;&ڶ$��W�]�����tY�_j"��� Z>%#m�:J��Ʌ�xp�1&^-�t:��kuR��7�WEל)o�B�T�
�g�O�`�>��N���^��}���l~鑽[K� �H���u�x�d����w����=���"���Ւ�f��7K�)��C��tJ?e~^�=�-���m��&>���bѫ+�NZ��J���;|z�&�h�t��db�6�3�};�5b3k�q���-��J�'�tG0f52��kr�Z|l�U��a�]��0/��(��'j|#���� 6WP%Oo\�b�G��^}����v��u�=����ziC�/۷�@c$0��ݓv�Ȕ��2<H(K�ڹ��G!1����%��ځȆ�]8u�f'U�7䅹��^���F�,��qi��5Ar#�I�ld=@\�guG�0�8�d����95PF� ߃��KM���P?�I��k#�be�
ȫ�sO��E��%�W	�����X��Y���;x��;�Й�� Qq_����k+����\����wI~1II֟�h;�������3��0�Ҙ�^����Q�G�E��lQ�]3�=/���̿L)�	Z"�5��_C����O%����A��JweD@K6C��&�B%�]��]��z}<|�Ww�ơ��z�����yG�������8�����{(�K}�_�����R�[���t9�����	&
~�q��8���Z�H�*Ԡ���N�M���i��G��X��*���s&�'�ՇGEv#o�^�+��uHMk�T Ǵ� �Q�"��蹩=5�-�gEr�p����?1��� �~��=w�����e��Ps!�M)>��h��;���町�h@iku/��j(��9?$�`/����m�u�g�ȫ�y��� �<���A���(�
<�T�a���^߲L��y��W�l�I�j��rD�ʉD�C�i� �tF�����%$I�H�̹HS�3�pq;��e'��������Ҝ���f\�e���o�ֲE�c�)�@#=y��MI&|�H��3���z��7p��t�ᨡ���]K�NWys��&��k8�<q��/��V�,��T��G	A��_��MW�׍�;Dȿށ�Gѐ����7}��(��w��EoJ����{76K�����7�X����G]��%�&V�����Y�nit�.g'����7������O%g�"�W�u!aҶۻ2�F�nB��0�L�^��)��u��J�
#$m�],�En�L���B��j �l��}D���W5��획 �%�w"1�����Jү��Ĳ��f�
�C���	PdLU�ƥ���"�Tg�qY3����K�6�A�9�x����e�e�<��QAw�����$�]k�/���4^%9D�,AZ��,�3�8�w}�L����EΖ�	�#88����x�R;Z����%�G����F��~��z�}�ͮg4��m>w�Q�J�D��9D�9pO�Ti�D�)4���u�"���0ac�����-��k\���� � �����2]������'�f�<��"L��\�/�E#N _�.5׬9� �m����pn��?�Ѭ@푌���?Z����\�V��.32\�s�Qq���:��/}�,^s�L����W�|����lx*L�ܚ��sR�l3����b�UΛ��g�O�,z�:����5Y"�
a�2[���r�BR�;W��Ŭ�Wԟ���/K���^���L�Xy��Y�kFy���f|����W�쵊@x� �f=#s��_�է�4K�b0� 5��@��˗�U�_R�%�?��uLk+���Xp��r���d��ݲk@���P��	��o�.}*���� �/��U�	�O����be*,�P��j�K����/��f��� �@ݍ�K	6A�?d���������7\���$���*!����ɪ��Uk��SC��p�,���rg{��[!�eu1}zC�g1�E<K��;k�?c��Uo���
�� ��e��/v$9#�/�ȱ}�t��'_�
S�������n#�O�3�#�{��E���F�@�Ǚ7�}!�eqQ��3�8nCK��\�dx�i�X�$�1�����<5�D�{�<a��
�>�d��ѐM���52���M-��N����<`q��q�$l�C����h�3�JF�u9��ik\��m�����0�{"�q��#g����oSÁ�E��u*�sl��&p�]���}}�V��1�)�D�t������Iɸ��6 �-[�mi�q���N?C�T�Ŝ��חi�Dn�@��v���3⋟��"���&k�d���t��Ym�]3�uM��6`J���c���=���`�M1�Z~���Lnp���`�)��M2����bh�ά)]c���۟��yo��A�Z�\3*��睞�ҿ|����^8��p���"'T��p���L��î�V|c��p�Ŀ��dU�*e&N���᮶��NR��=���:����h��]���j�J��$���+,,���kaÆ�7�	��R�ى�ۓ�ڼ�L����������%�%Yd�n�,	8�3���E�����Ȋ\�\ Ir�.GI���*s�v�Ǖ�o��ߎ�M�]�~�Nn_H����{������D!%��I (O���-Sk�����z�.��<��q���.`�,d��̀A�N��ɕ�fm�EZ�q���J3#7v��&5����J^�_�Om_j�\��i�JK��pwR�e��u�s�'����S���s�լo�����<���B�Q[K��=�G�\����M�?	�b�m)�������e������l�ګ �'���4y='��-���{YyA�,�ı��t�r"l�+d����?T]]�7��v��M��Q��15t|,�t;x����#sO�Յ �����}3�y:;�D4��<���l��0���>���k|z;������ӓ�B]%�t�|��Hr$��jT���$�� � д����0�p6���|��0q񪀎g�X�rv_����f>N���J�\Hj̓����Ir�D��(U2�h_���F���3��]�g9���N� ��=�.��,�V<!�i��W�������nVDVo��*P�+_	e�$Ƭ&��(��*8p�Nz�o�Ǚ�G����e���B�򴸋[��Q*�. X2���t��:	�$%NlKFSZ�f�&N�ϖ�[��lu��S�YӜo���⥩WwL�~��J�w� D���K:]d�ݻ��؈Tk�q[#P��zGc�]�+��K�
W*�����ng���Y���mIa2���s����X)<2NFa��������j�Yv.��2�J���xah!b|m��jl�Ccm]��͙�#�୳@a�9K2�u!O ~����F3��ݗx�p>I\J���#a�Ù}<��	�ԁ��/�����ŀ+&���8vEy��}�����
����o��VA����ۃ��ۀ�,<wA�K��/A.�R�{qCJ���ÿ��H0��.^��H�S:��%,R��M��J���}ճa�F��3БF/a	5285J����ՐD�Y`-��p�e��WH��ň*e�a�%���'�v E����'��>����S��v2_�K1��E~Z����dUT�.-n�O��+����d�W���!l@���z��a���јǼ��d��<
]I���%�\IN�9����:���6��0X���01�y�ɍ&r�KT���P�"͎���~�~{��aHY�g���#ؗ�c^hSӟ���"~�3��òz Ӧ�����fKnϮ��+l+�I<���	8��
+����d8[�.\���V�9�^�1�A12X��o���K�Z|~�12R�l*������?�+�a}!\�R_�:����Ի[�K�Zb�(���6��Q@wĆ����Q��:ݟT�����ej����ӥ$)��c�SϘ�������vS�٤��!5ޏ�I���lE7�TkH�@0���8E^��1�h1�\��λ��@��kJ��hl���Z"���1ж��e�u�������i�z���⮦ c�)�gh6�������7��o��#�!�����)R��k��Ԯ�o�J��l�/��� {�:۾5g~��K���� ��l�F[�
/��Æ%Bi��|���*h���5�ҙs�Ӟ*{�E��W����P�W-}Ľ��Kz��@�|`�GL6%�,��-H��R���l��6�8��׽�߸2)}�#m�ѷ���,��Qz��F,레Iڑ��OI�@�V��d5�	�s*�6�{�|�i����ST�k�;�t'�$�n���m*��%�3Jr+�B�BA ���M�{
.E�ά�z("� ބU-w6���"F�s6^�_��m!���Ȉ59|EJ�����XSt|��xa+c'e�P�.r44��Լ��_Ҳ����7�
�p��l�l"מ�ݴ�l�ΦH0�3�T�W�0��+Ҥi60@j�#N��Y<�`��K^4�4�F�zv�կ�5H�h��<� �ow�i��S���PI��S���2��c�q�N
`�z�<�}���dJ���:4}E1qQB�Z�"�e+�����f� WF\{��L�J��5G�m���hJ8����[ �o�B�������+	n3�&6_�\%�zw�!�~�5�kjpV���-Ǣ¸g�ulv�/��f�+�lF��T���X��?�[$Hd���eKײ�1+�4D@��fT��$g�<d�(�2�y
Z1d�@���%�
8	#�X��yG!&8�ia��9<��}��M�3\����WW�o�Z�uK^�3�p����+���*><��Y���.F�;�}!��R��2֨�Hp�MN������|�-�k�w0�K���?9T����ijj��3���oj1-b��+a��.��*�:W�T���i�-���O����E�x9!|y=��Y>�FZϛ�R(I`���-�b%�ΧΣ�/��G��8YS�h�!u.�b�m-N�M��1%���0��
Ne�D�ٿ[:W��_������Z[������qf1�������w.ߘ�@& 
��J���cI���sTr�,��R���$�`�M�('*y+�XVC�*�����Bԭ���(�ר�̙�,��-:ȓ	�|� ^�.z�V^�/� /�I�:�����$�g3����tcI^�,���EYX�j���7 �F;=S��T���]Y��X,2�`T����-DBJ49t-���R�^�d�	�mŕ�~�ʕh��}2��R�3��"�#1�BC�
�Vg%%�eۺ]��i-���	��@���ߪ�<��*�|%`hS�9�\	��'�Q���h�$T�ו�Y5=���P�ĵ�:8m�|l���:x���������T����â[�߁����h)�$��t�2hSc��ː
�Y�,_<�:�wvw1���y��4��B�A>��l���Ǥ�]ұ:N|� �Q��d�JI/gw�Q'�n�s} ���o���Q�\����h@��k7��P��1_ �/`8f��@B~1�I9����tT^��o���
�%f������F��x�h'���ӣ�z5ĈTqU/CN<w M����v�@��9�T�����:��n�}�n��ժQ;�iJ�]��]2�R�VS�a�KG��&�K!�Cw	=$�k�z�_��Pb�k�����sȧ��C�`P.6ÏB�ѐoSU<���z1����ؖ&�"�M`Is�z�_M6�����Y99|��-��A��j�R9%��j��5u3iF d�U~�S��P�ǟ~�r�$��4�w8[������W�~b�;F�U�,�֊R{{k��VQ��ժ�Ѧjת������ﯓ?N��}�����u�s�wg�A�cl��/%���-��`��z|�4��׊uJΛ�#5�������TB[�JGP��X��\���v���=�V��">�s�Y 8�<W��[Wݩ��~1Z ��E��!Y�g�eӄ~��s^}�ޭ[�57Q���g�^Aɛ%�b�R��H���0U	BK���M�Ӆ���	��c}��&|c������C[v>-��8��Ze�o�0�@On��)��3�#N�e���"q'F�i����ܨ�u��5�����nO�n�0�+��у��a
2�긧7���J�5T��A�W���	�M��(���Y�.&�������������'%o�B-�66�I�1�*z\�s��`���77��>ۭ���/���ʆn�w��?x�û��՚�`���)�UB���Aj<��|���%A:���񪍞�� ��].��$2c�[��Qk�Ģ�c��T�x��.�>eMi;���ݥ�E��N��?���8_����z�gf-;,"�ɷX05��9O�,�&dȭ����NP\q�P<��:��6ZTx����$RR�noV:v;���uKZ3���<�s(��E%~��� ����������J-*����e��x�&h#�O�~0�P����슢�D�2.�au�ČBUET׭!9�����ھ��ſ���qn�z)��'�sKQO-��>���e+��,G�*���%���(?�?xM�9��}�����z0K��(}�ڲ��V���e��>�s�2<�Й�ܛbf>���"��� ���t�Q�M�_e���^o��U�����@&��RSaػ?O:ib�Y5� 4ċ/���T:/ȃ	�"	Z0�<w|���?�c���ș�ҩg�q�j���9T���U{_bB��)�*맫�M��O�ZEІ��o�D`�l{���q���n���TIog:|~�9�P��\S!bNeں,�)���ћ�䞑p$�:��{ x����>NNHt��8>�p1E$�Vz,��X�����j��f���xY�}m ����c���.��u�]��ߋk�f,�f]�_>	ħK�D��t�@��Nk#��{KoC�U��A�i��1X�iR�4�>{�gH�f+6:�kj;�"�7�Lk�d m�S2�N��D���#�Q�S�X�jWA����0@���=��{�y�PI���C7�wZe4B DD��B}�	�$u�3;�s�F��HM¬#	�����T�����������3�]N-���_zFx�IC)A&侾h���u2u�nm��
s>r�;A�O��m�5�C��>Z	Bn�������'Z��	������$�O?E���5�����e0�-��c'�ڃ���t�&Y��=;(B@�Bj#^�:��	���ު�/�NM��E�Tf3���|�UI�}�7��H[V0q���!��E�A�7��P<�����E�p���Ȉ��(��]�i<�;r2��W�l���dH������n<oG���v�&��%i	��r�i�f\�v.�Y6њ�4�k��S+MH}踶�-�1������Yڐ���vG��8�BG\l���|I��YuKs)"��O[�:cӔ/�vg�Lu�u[�z��DG��8��uۼ��l���6/`�K�_5����ܼ�����d�?�sʙ��X)̚�`2�GR)�dX�%�u�Y�V���+|+5�HL��]8�6��F)��������T���C�.L�7ɷe�Ō�͛�oR��wt�n�ّ
��TmJSq9+�9o���b�"$����ھ�G�O�_�ga �щ�-ݍ2[�W�L-�҉N/KĕP���%H���D^m��C�~���0�Z�a˸���Wf�Zj�v����ꀽ(e�;\֡������2>�n^6�Ƒ�H�л]�S��qF�O�^�}{��rŚ���預��BC8E_�8%������/s��j��5�#���_��7��GM��($<|xx�ܞ���Po�ʆ�4kI�Ԙ&��A[����\~�B3.�CWv���X�^kCI�E�)�Y��>�������n)���2~��s����Ε�6�����z�K��U�M�-���`��o�h�l�@!O�Γ���Sy�o��w�Ő��ݰrs���$������O�Y"C�L�ĕ�N�����te�we����+��&Z��\$�;82$<ǅ �A��ԝgZ���9���@
 nzڧ���k{f2��
!�����i�f8���޴ɋ���3ӣ� =y����&�/l {p�).�6Iy��:�֙�{�X��=z��׀��GN��EL�x~s���Tw��Əd&h3����*M�QD��X��!�I� S/�;�I]�0�Á����]��UC=L��x�A~co�&bb����u��A(g-�b9p�Ao�cM��8��;���o��[���b��np��4�d�N��2sZb������X�p�,ʫ������|�%!���Á$��"�eO˽��}���n%2�Q(]>S	��F�P����o�(�Bj (���n�6��={��P���n%q?�Y��4蝹���K�M�ѹk�+W4(�i���3566ub�g:$�?v�*��S ��oQi8�w76��\����yD�
�jO'�8��K(�trSF��/�=��?�=������3��S��噅�s.MK��wv葷��̳%�.z��I�/c)i1P�#� ��Z�!
�8�[�Fo]�N0xp_{wgT=��@���?t��!f.أ���Ed���V�/���E#w3�Sokmv��^w,�F+Nx�X��»P�S�K�^�:���o^�KNg���F&��:{z��.7���X/ې�����
��<�4 �T��{i
�	w���^��
�".�$M��%�V7��p)XS��+�D�
A��o�\�gx �D���w�iyqJ4�����bǄB>X��-Eݹ��$�"I*�mFk#."
o�v�~ʮ��*o�~��!چ��dVZ5�Z�p�u0��cGu#��Li�ӹhp֜Ϻ�N���Ê�Ev-�L��JII���Y�l=5F �.��6ý�2'��.:R$!��E�y��%y)b}�%[�= "�P�@�G�>���j<�Qm���a��d	��T�w]�{ٛl�侤p��5�.u55�mu�q���s�٬��U?8Rd�1E2L��.Ŗ.�(��l$ �����Z>�Qof"}ҝwc	��Վ@�4��p���t��CCS���y�2��:���U�,�s�ɴ��Ϟ3�Bk�68m;Z�4,�<���#������������\X��
7=��Џ��P:��E����W2�A"bď�=?h-��uΈ���>�J/�!�L�Pp�s�7��]�3
Iy��|�6��	 brA\��0���xNUQ�L.L�������q�@𮉬����D�y��o�)�FY�Ί-�����q�=��и�ԧ.#��&��K�ڐM��G�K�z@ #�?��-��d)%��|.H5����v�AD������NS��2�s�'yW�A#v~�'p�t����i9��/񫜡(�՟�1��q��^���R�H��
���%p���E�3>jM�}���X�)���o��WY�r���#W���_���h?�|�f�����f���,���t�%I))g����aE��
�W2�L}`n~src�\�f�X��H�i`����Wi�l�[?>6ߥb��XnW�*�8��G̎��C��V=/9��BKB�w�n+�|��d���R(�{+MV��X��B��7c3R�H��"�DCg$Y(���_S��5An��ҩ��$���5EKg?S|���5	1��W��K�ȓ�s���˧W��z?'
��
{2*'�^V�?�O��b2�ԓ�HM��i���ի;�u7N
4X��x���u_^5�߰�f�T&��UE�.�h��vMw��U�ˌ��P���dql>X��&V���7g�/U��������
U!��Y��;+�_|@��H�����6_B����Ʀ���Y�)m>jBa0Ù �����k�k����	�8��J��0J�aaq������Ǉ�V�'�g�ƶ�|��S�>�M��t�"�/��o�77w�3Q@~���f�Wx�������42�t1������{w6jj����p�'�$q��$�(P�ߍ\ٓ���9�[�B�㫴q�5���KT໾{BaĽ�D�'�t�6q�9謳4��
��PL/^�x|sC5}>;/k<9��R��'�k��!��L�4�tE�;��T�����0X�E�-Nh�i�]Ğ�/�z>�ONR��,�r^=%��0�x�w�Z��0�u���[r�/Pɾ�p����Ȟ5YA����{��hj��./���*B ��cK\�ձx�f�L�����������{;�>��\ �oC���'\�g���oS*��z��w9gPD!` 6:�kZ������,�����Y��W�~�Y�oR��o�[h��SB��bk�� �)�����n=�ŵ��y�@z9�x:�N�}�f��^6��t���맦�%>z"{�9��j�+���֏ �,��Z\yP�d=�|I<*A��J!��6c�������Rq�H�s���z�k��y����rqb4!y�?2�"�A�� G�4�3-��^�qX�X�mA��9�d롪�O9Sx�����h�.���q��c;@C}я���|�:�/�ו��Z{��I��vd����ٽ��Rt� @V���"U�Yg~B
ƙ�+ej�4(��v�����hE�g��@��N�hߜ84IJ٦�(˃F������g3�.�:Q���83���s �tY����*/� ����+vd+�5�9,��_��Q�[2�-bӤv�|d,!����������y�Ư�)�)�1~��^�{Z��N��$�Ͼ�����F��^ҹ`�g�f����������l}f+����e<:]�}�4�;�T��Pǔ�I[������C{�G7'i|���_�ZV���r�vw��Jm��'���P�/�l'�Yb���_���:'��k���j�^|'����~�a4���B��"�T�����!�5���2F�'��x'L,86A/M�s:@�*N�����"f8�[	Uc6��t�+v6|_C'W"��u$`zI��[R�Hr 8����=s�@��~����!s�>��-sO}N�q���G�MFe�~Pjt������*�l���M��6��@g:d����&g;�r���rІ�yozt�r�	V&��&i�N1�܀���m����6�&�J�:��f0zx���Z?��S�p�B��L'2�:v���B�v׭tI��L6w���Ҭ�(nD/,�9�t������r���]�f�9��5m}�N����.�g�o�O��_0^ۨDS�>]tGgo7b�4ߖA_L̸���:�3����(f��͐�vuʅ�9|�?Grt�d˟� ��%T9A�U�Ŭ�+=���OƓ�{]_�}�����*������^�zҌ�zʏ�n�/0�T�OY|^Zz86�4%&�
��t�*��8q���xƛ/66��YZFx��č������Y���ճ5{
�pf�?�1��N�T�RM���H���Y��?�+X���m�����rH��I@�� 2Aa]�;��o�zF%�����OJ���ʽ�J�I`�}`ʈ�-3t@���5� O����ǈk\��F�0�$�f7��)����T�ւ�1�2+ң79f['���߅[*4f�D���_Ips����V���:���8N����7�/G�*��;��D\{i��'���N7���`� ��NL��ھ����R��P�~8@(Z��!�Ќ�ӑ�폌����4b:��jZ��j��jP}Llq����PO��2'��#��d
Z��(6����/0��.O04J�ԫ@k nE�[�eIvD�����B��Qr��I��<��+�V��U�n�	G����[�����*�Ggg14�߼l
�!�+��&Z�/���b���L��|+��T�T5���{�S��sn#c>�\擢�t�z�FCY2����GfE��S�`@�`��9O��6jq�n[�� IQ8�k���.�q*+EǾ���@!AkŮذB�_�	+�� � �=�tq�XVֻG��(?�*om}���ՠR}G�ڎ8���Q2�C4<��2M�m���5��R�\|���y�$�y��!(g��{(,������"I����ն��֤J���O��6���v-��(?#IU��V!Fy�@	�(�i�V��3 +�Z$j)����:.�Ҳ ��.X��Ŧ�3���b��|X�cw�O9{Y�[99��5Xq��F�v�;o��>��fbM��]Bx�)�,�� �:���6�Z��u̷L_,�㗭�tN3j�U2-���y&����څ$�d���ȕ/B�>V�p�yN���~��$�v�V۱g�@��@H�Ď�Vwn�� A"��[����&�ӏ�Φ�M�NwCTv�v��Rx|���r�[6G d!��C��!:ۂ� %����~5��~3 ����\��$��yJ3�I�dv�{��m���ZWu�6����ҫ�� �2�2�a��ߝ7�����~��Q�b�@h\�Xu��y����ˇ0͂ji���Z�����h�5V<�ɑ_�wx�3���F!�b)�o��`a3������Q?�P�7�%���]�:&�K��y�����\�q�irp�A��t�m�,�;�t�d�Zbr0�G��jy���+g��cZB9oĈ3�?4BB����������;:�tٻсvlw�T �y�k�\�$�;��c�|�N#Wh�~��g͗L*Z΄�Ɋh|�A�cS5i���.�x���2=Kk�� ^��.N0�2����B!	��,�y�F����N���I̗̻b�L�oh
��H1aϖ������.�Ag��1�і
�9���_��y�X�`��5&�Vz�yѶI���f���*��n5�	Jh��]X_V[P5l��$5�Ĺ� ���R��a��b1��n�BM�Q��j�/?�R�"���FU��S���7��(�V!7%,��{R�d"��^��!	���v%�{�#BaX,v�����/G���k����"i*F蒆Ÿ���H���g�x�o<�3�.�9��~��
�o�T�4����y��5�K������ ����ҭ����ї|p)N���u\�P�����	 �I.ZA������2b+H���YEf�xX6�)��Ge�D����}:��1uJ�`F�_|���V�d:ʈ���+�Н)�� ~����r�����#
91m�CAN�)��-QU���3�ʥ�dǓ6�$¿�s�>�Lo^��,F�����c�"o���D�^Yh�����
�^Ho���nI�-��'��MDAk��8�_Iv�v��?�\}�!:ؓ%Gȭ�ǫ���AJ�}�t�E�[��V������3�\(�rPZ.0vZBàFV��G�:Nҿ�S�Ţ��  �%t����pҝd|��w����kdo]\�7�[��T�q�`3$�g�����˗$�����5'����J�E������xJ׉F��������s����C�v�n�P�V�h�ܕ��KB�I���ң݅���/��~C�sΟ����f'�Y�[A���e��æ�1玹*=|��]x
�y�-��9�x%�js����|�-v�/B�g2��ɳy<66�Q=���[@=@R 0l�e25��{#�b��~}�O���q�ܙ���]���������ݎY��o��4��U�C�Q�����A<���O�F�1J�������-dD��l2G�́�1[�;�Pm��(��4g�7{
��'��li�c���̿�c1��.�J���8��8;���H�a�:7��3��@ X's�X]��wk-wl+3$/ �'v��Y7O|(��C< 1�"�4��.�$�!*|�."�������I���RW��ݻfd̀D���Tؿd7x[m4uCG����������b#�K�d+�m���{EXl�j��>M�����1��W���[rЬ�Џ��G�t�v�-��Ą��2T��K�P���]���Z�pnmu���@�/[��>Mt��'�����!����u�*o�
h��A�S>�>�讻�;wj������:,�0�O��|��b]Ȫ���hx�2�B�CHԤ2V�h�[�lc��X�`8/K5ģ�NudOZZ���6�h�*�vk���ih��rgbfl�sm�}Ԣ��{>���g@��^��μ�o��Q���SHRi��ra�C���U���&�,�G��L�͙������P��Z)A�͹�J��}��6^A������9��1f����G��b�E�D��Y��)��[���"�^�2A��y�#�d>����t�켵#A���ϳ�y{nZ�6��j�z��2����TPD������V�3C��X��2��6i2.�+St��
fhr�R|rpsSP-��G�	H-&d��_�G�
?}逾n�f�l����/l�@X�Ԃ����`Y���V[����P��vht���߿��zÌΥ����W��U�3J�ss�ߥ�߸A8�XI�D,�^������ q�����[��e\p�O�	���V�[�;o
��a��z��l�oKlG��d����r/v�F��E4:^��#j��թXH�1�z�Y���%�����_�d#J7����Pژqr$�+���K�����c/L!^�q3��#ZBZ���q����%�ډ��
�E�d�}�kؤ�o����F�cM�Sm��z�5�%�wVA�B�Rp�?�8FZ��@�;�� \Ȱ��ϗ�W4�:�č��Q����r���u�������m�������:��j.�#+�l[���ѱtS�(\��Ұ��#���ܒ�U�}�άE�f���x�0r_�H=W�5*3t�y+��������b�zGs�V	#�N���JL�;��:?�?t�ʕm?|}�)u�޸�V�~{�a��:�\7�G۫��/P������<ܦ���,����:�$�q����JL=ސ�"e���U꼒���)��uv����:��4��p��0��T)�W���;�26��䘁����֞ך��RF��J`��w���X��'77f,@]͵#����6�E.j�Y�a	G�."������y'�;8�����ǉ���/�v!����j���A�؃�$1߿Y�]�vg�$fӒ� ��fiU��<�����[�wC�Tqnݺ����n�im�u�L?��d9�`��הE�^�^��Z�v��X�����B��X��A�fpM'�J���B��oST�˾;�����?���F]Z�(�F�;��i	�ߺ�9�mu�f0�ھ���� c��Gb%ui#�GX�ר �p��Uࠟ�;�h�ɪ/^���N~��E�^��'�µ(������eS"�V�׳%L���ԓW}�\����B�<Ķ�&,������� ������ײ�p�^w��I�Į���5�!�`��˕�6��j�Z�I�4�3������f*muj��Ş�9#ƏÕ@rU���Ƀd ���r7����ՌA��h�TTU�?�e�:?4��O�b�t�˞�����U��uQKB����tt<
X$�w�ɟ�� ���v��+݇�2g�w�'l��Y, �mD�����=���EB95�{Q�c�~�|>�������$|8���Eޢ�� �ut��h��oU�C!�˙�<	j�O־C_� �����4v�w���BH���r�ݨ�j���v�'�B\�<��������)�;yU�2��M��z� �/��ß>smx�ǦlP��ې�?l��I�w��F�d`�S2���$�i���~X�xQ鞦9দ����ǘ����y���۶�(��f ��#��F�(���e�W�~<L`ՅK��C��#�z)?��[ͬ ą�/���K����hP�ޱ�����RVy�̢G�w�>Jk��4������! �O_K�fK�I��2O
K)5���`?OMQ�`&,�X��� �ȗh���뭤�r�v+���В���/�8@����^Ծ{Rѡ�MV*-�1̆�	��I�3�ϟ?�"܉��D��5��F�T���,��y'��%�x��Ǧ�OɊS%Z-�F��~P_{�����ӣ'm���t��S�ޘ��7	׊@(�4 4cc���CҞM��Q��c�T���Xo�
����~�^��̏0Q�qd�Bw��y�uU:�h��`$�W��-Dp���[	R
<�Q�$����#����St�L���n&�tr)>&� F=�ɒ�_宸����Tj��B"C?KS]�2�����:@������Ǯ�fG+�k%����и��;vz�*�����{�=�AV�'��m��Q�9$��Liy�Jiǅwӯm��Z\5�D��̪�QNl��U����F����.q���0
e��S��.}��s/S��b�3ma��Ĉ%�4X	3���O�@Ee$m���<�0Q��CŜ�7�~;-�S#i��p.H�s[��;/]MF�u����H�gO
]8�W#p�w���, �Kw*� ��C��s�4�_�H7y�m+f!`�N��1z��jqAFzL�uLW=K�������:wrfQ��� Un4����R����]�<#r{�Z ��#ݤ���	�޴dn�a�!�'Ps��\��U���1�a����(��b ��P�H-}pfղ�	/��f�.�9lO�(���BNk�3�&
�p�l=g*�<�y����=T2]������^hF�V�׸��oi;S�o���4^I.�b�{d�Ł�u'B��Q���<X�+f����4VXC��.���<��1&��]�٨���V`m�VG��<DB���֥˦|-������X���mK�hį�euuKR.Z�k��i�ѻ��}����}�3R�߬-�M�6�>�H:(H���i������%z%����_�Z9Ï�ͬe���)��H=�^X�Yi�{9�)����xJ~yn�Q7ם���C{�\��Z�7�t�"���ZDdm�	MV�$��}S�"��)�˨ӗw�_���a�#@I��z�ao.�9��Y�lC��>��%�w���Q]�-p�[�-����oq��d�&���t�-i@�[��|I���P�Ċ�?�ݺ�e�J�0<�D������֋��'3�߹�F1���Wv�d?j�s-Oj�hU�J�ܲ� BG�6���mmt���������xN�j� �3������B���r]�o%�(�Ӓ_��[h[�����RRB������Q��.�֙�JSq`
JQ(���?G�t�T���G?c%�gM�4��T͑F��˽�����ҁ��wj,Wz�};[�Vr�5�0W��e��Lg -Xǥɮ�,�#��~ ��>�7�����R�x���?Եm6���WK��dԆ,��>�s�@F�JDR}��Io|4�}��Ѓ��BȜ��&�g���5U�<��!Nٮ�豍9F�"֪.��7����Ϟ33,��x��A�K�qu~�û� 7[
^��`���VT�ƅdW�H�!���e���J�M���h�"ͼ�Ÿme�˘"�1|Yܻ�G5�ƣ�đ0�]Pdh�hS��G/�M1�h��a6�~Tc˯Z�iUէ�{|v�2�
~A$���������
�=.�XF�Z��8G��?T�Vxܺ���}W	ժ�3ץ�d�>?9�ֻ�����8^�|z��G��I5IJ�(Ij�o\YI����@F;�V]�I�<�I�49�8��:������UF=،�M�z��8i<�	F��˷�*Q!8��*h�Y�5d�����;W��E,+
��G�g�y��V���{���D,�Q�ڂ�QN�1��r��N]�ݯ����O/��n���p��эCF�:���R�E�Xc{�룾�$�m�x� ���-�r����J�Z�|����i*J}o��K�g�wv�V�d]^/v�c�vp����d}�����ϷS�:)�M���he������B�"L���8�u�d��m��\�t��� mL̬����}��鱋|��S���l�t�P��EՙAw��5,m���C�/x��!6��4`�Dm_�@!C�BG�֋o7�L���3N�jު��2]�ܱi�𸽾O�\��`T�t����"5)��L��+��%�ؐ�xϣ�R�q�wn1_�Sš
f��]���܂�r���Y�c]}��s������à��+p���Z�H��$�ӎq��P�p?�A%"�"���y�bb�S�k����ٟ<P�	,ֆ���$��0����Ŝ�V���u��w���`�8���v`l�Q��l ��:�C3�↞B�e;%LYoT\����YL԰~i�6h
��bo�/��S�t�Gq�Y'Z�|�CX/-Z�ϩ��B��i��6�xX�-$)%e.+��;���r�M�#�.�UJ���e$�����U�b{9p�Tp�#,�6�����E�l*���jZ�j��߹�غo��?M�G�>���7ۋK?o�����&%.S&Ռ�7�H��HB�Ϻ$^p2~P�j���\�V�3R)�B]e#kb:�֬@�`�,�٬Dw��9w�/�fL9��b�Ƭ��ׂo��"Jf��'��F5鳚YU�9Jl���K#����U��b?��V�f;&�,�!�=9����c���x&EF�����6
�o�s/A��ThJ�#|��9硩�DW��5�D&�1#�y���ĎJ���*ʂu�i\��]��*�����jPe Gά�I&�K�w�4�7ݓF�%	�,!	����Q9��s�{ů���ئ��-���������"��G?�$++Xrm
��E�Qg�g,�^B�,y�q�f"j��<j��⺽W=�R��%�;��n���B�&b�V�g�m�>�hFe�t��)C*(���S��>�:�'�����j�1�?�DQ�y���n�I�3Ӭ|��@�0�"qO6]�n��	-����۲	
�-���+��`�P�����n�Ċ����Z'��O��E|R1�/��?�,H��6ey��b�E�Y��Q�B*v,����D ۉ�R�2d�pѧ�:��d+.��"=zm����9����T���b݌���WU�S(���b��O�H�y_��;��=$x!"f�+az+�3��~UI�ߵ�S6III?%K}���:���5�E^	���W{{�}�����~�q�)Չ?g��&CK��������p5�Ҫ9rt�D��o ���9���Y�����v8r�"����H5�t߉�@0�m��R�zwV%n ��+Dn���~�i���I� +�2Тe�p媹HKL}<��ż�mZBl����"c��N'>?��WC�anItJw�rym��9�SI����?x�e5k(���}�����M3��N��}ǥk�4�X�
w[����ϋ��jw�{
�+
>��>�
��#���a.2�W��l��ۏ���Ǥ���
�R�h<���4�?�����z7��̍�*B����v�v3�u�$����.��Pݔlh�ލ-��W�$-�~�6b���Ƙ�r�9���t?�S`�(η.�PW⭴�w�(L��>.i�������������#k�wA���d���>�~���1�)[Ƀ�=���ᑡ�3B�1�jq͑�Uf������$��' �I:�9�sl2�w�&���
��y^�p�DM�o���(3qn�J��r��:v1n��R����?{�bH��ΰ{i7��#)ʉMtU,�����6��@�|����}�Il-2]�5p���+Bx�� �I�5�v⫂�E���xiV�"_K9q�AI�9�����G^h�\�|�;`�~Ǿ�+>ɟl�ܰ����C�m��>%�~P6���b��Y���_�]�ӈh��
�+d��>�H�i�/GW�����Q�^m�Kh��<J=��G\?�(��-��AS4��Gc����;-�=��V�j�f������\7�^�3� 6�O��5��~e1��%3�K�]��Iҡ�U�2���Id4䃾<$���d�>9��YW��z`hsD��G#'+Vـ!�9�~򡽃�3��JD�䋤�IJ�Y��� 0'o�gHi��j2�k��p�xhN�k'AG���Xze��F#h'amf���l*=)zL]"�y���x;��tfD�;�,Wg�y�cS���fJ�󶴸��k������J��$�Ă���XW�1�q��Ze�n��/��'�����I�qR���K�(�J}S_�/�����,b\��S�c@=57G&gG�l�Ƅ�wG��S��O����83�~x+�؏�ҧ�ǽ����W���1����6'3������l+��4X��^b�n�<j
�#s�@mџ+�p�h9X�	��4I|n���X�5�e�Uc@����+�A5�XwiI�S2��tS4Ȏ�n^�h_��ĉ���s��O�cZJ�,��3� ���T+�Ќ�B��3���?ٍ��E�K'����Fh���UpN�{E�C�SBII)N���_{���rkk�"����άk���[�i#|9b�;|�)��O����n?�Ն��5=����>?4/`�	,��h��=������j�O"�d��:�:*^�!�Y���s9?��!�(��_#���������.����Η���ɇ��4/���{]$t�}xxH���V4�, He&=ܓO�0X���<aH#�/�׵�tѥ
)����	���b���e)�
1}q	��(]:��w���Ƣ��)#ZC8?7��*��
��ɢ����?�<	����P�[�+�_���x�Y|:N)���)�	�Z���(��z&�DB d��m:�����(4��K������ƽ��ZTB|6pjo�0\�by��EZI���w�h��͉�Ue,��Y��!
��$�U� � [l�5�`�3�W���1��btTO�� JiwbW���b��J�7C�.�Zt�S�tX�H��%Nڳk�I@V<ԯٸ�J7D�z&�Si<�x����Z��+ݒ*� �+�wV��̐��s�yh��e�����S��?���SWU�8N���K#X�.�SS��0��N2��>�%*�������ښe���Fy$�S ��ߣKOX�$C��+�
�&!�w\r�����d~��1M}w�`��'G�5���h�J2Gb��"~���!Q�`��V���U�����1�pe�2��E{���,ݒ�ȍ6Sk�����!�����5��×��)�3���!�V�/�Y�Z��VWcl(ީ���'6�c' ���Β��}��M��6m�a_����S	�z)(x�G.װh�f�5)��O��s;	�����O^xN�L{tr�@dAj��&�K�Զ�"hr��Z��,?85E��"�>x���J���������!>�]�_�w ���R����\�T�I�iq�%��3}�6(��_��;b9���Wf@SÓ��X�.��� E�
tj���,F����
�6ukYq٩H���$%Ł�1z���O��wU�dSy����#]�����r%���R�/u�qO���d�f#�r�{8�},�������H��<���(���{�x�=6��Ge?�?�#��2\�"He�R7zqO/<��ɂ�TȈP͝�E靌e>RAp�p�}���C��U}��Bi�?ku��dR���� S8)�f�PN}ݢ׵J/���qMG����;v�?}����kT	N6Dױ��!,f�'�w [��bp�2ڃ� V�_Ts���x�\l�Ϻh��(��_Jw|L���5�� ��̐�:���p]Ũ���?���#��Xj�_.?&�6_�.�)��ذ%�.���K�о��Z��~n�^%�y�l+L�Yl"��
�t��罹e�t�7�M��|��Eks~�Nvp�"8���&���D�=9���{de���1��W�Y�1`�b�#���<���<|��3m�pxM���6��Ӌ`��q�ٳd���������.m�r�f�(9�ڱ�ȼ��zx�a	[HI�۩��5�dh`>��!]� \>/�V
�=M���r��)�P�"	_��x��!����$q�F�{0�/WG!F����L��`< r\1��n�{�P�QK���NY_�[�i�_�##?�U�uvw�����q R"�Ij�"�����I�W�[3PX��oNݍ�{pG��Q^�����P .�~�/C]���є���4����#����L���$��ַ�(&���@��������+4mS���p��]�yDR��᪂d��������Q�֬�!���&�|��D�g4\��������F���hA��h!z�ޣAD�`�g�Q3JD2JD�5�y&o��Z��Y��{������s�����~3�T�^~ۧOy���L�6'�dB*9m�螎W�O��S��J����_
�a߱p��ZB�Gzv>�"��1gk��x����9��p��S�t���3�z�2�&�����$~����},����4�~Y�}|43��QbK���!�0M��{a���O���Q,�]5�׈w�e!�Ky�$o�G���c���YQ�y�*w3�R�g��y���5H�0UC���spo���
>[W)�2t\'4d�[ؾ�Ӧ6���5҉�@��2�#���q��3^�ɬԭ���a/�B>�Fd<�ir*$�^Lk�E�Ԓ5٢}�i�4]�;�������Ә�~��(�X5�ɽ�~&�L-���opa�_�'9��>7a���^,tI|��N�q,b�׌̯�o��_����k�18ǻ͎��P`P��*Z�
���%�Bǡ�T@]a��n -J��)&��Y��)k�\Tn��$�ߨ@��Ȭ�/P�����*��I";�� �s��>.��T�& ظ�<�-��]OŴ	O[��fB~4ZoHB��F�JYvw,%�{@�ϳk5̴�M^I3j���W�������5쥡�@�I� bt=��\[�8�j*�YD�1]ӬQx�L�3�	��:`Ou'@ڲo��`	N�w4�_��س3b(�,s�Ux+=�
	�����$�J���I8�~���H����җ�TՔQ���́�ʩ
�A"�K��Hr{�xM�j�v�ػ�uak�C'��ݷY�|7��qwC�2?>[�΂����K�T�۸ֺcam,�@��WY�YF����<�����4V�?!%~��6ꦝ�W�� �y��73&� uO��	���5�������G��7�S6)j̣f�x	��2\4L݅|�~�A�u9*���^��3��߮T�8j���=�z5�\�#�kz��>O�ۙ��h��x�JN�w�}&�1ẇI�^:?'E�8K�� ���$A\Z��4*#Rvv���]5;EZ�q���������6v}Ҵ��]�v��x%mg���I�!���O����������������f�0~Z�E5��j�Lb$��,��-��v]��c�C1�����oz�ݟ��.�#zW��Ti�T���I\��Y�N��3(�R���\!
���P>q#mL!��jN�;����\�%�R��4�2�,�9^���m�O*ҁ��O����Ҍ�J(��P��+֩ubDBa͜j23^2�u��܎�d� �.9���Ip�����qe�
���Xs�-kU�d"�r\�|��WK���(qL@�4�����U" r�vp~/�,�)������4��	V�6�зŀ+�ן��xj�<|�70pOġ����p�tm#J�k�z�'C�=N��$�Ԩi7/^�_����_�|1��M�\Ϻ��~��6y���:<��1�2�D��;��!p���Y~>�	ү�)>I�
J�Q�XZ^V�sF�zN���N����E�b�W�d?�8�9�[��Lm)��?~���BM�g/L3ui����&��y
�xH%?_���[z*rb�s���.��y��x��m�i~�=��s��N{ ���{~��<z!��������v�Fz��F���f�����n�����]�I|�rm��]���ֆ�u��;m*|{Z�n�X���ޑ:N�g�]Z0��\�����_+5S�k�ë�*���
4�ݫ��7[*��3{o_<�zQ��o�;��Ե�E i�3�ʸ�Z��r	�e+鍴�W��G�wa�pk�����Y�p"Ѯ0"��Xˮi�m�i�EKm�a����(��̷�'�?�d��	���zu.��wE;~���*n�q7u���Ӷe�??O�E���y�Lb�ʣ�VIo�G�B�D�q^���NK�)Z�4O�n9@au�X�C��ԁd��/wv�ⲕ����(k0ِGw�y|����Z�`���s�@��y��#Ҁ�2��c����ѥ�	OMI�8Ä��w��c�z��"�X�rW���X��^�i��?K%_$��||Kװ�7�Y=Ѕ�(�rq�Ϊ�V�.������	���:`qб�U�[ ~b�M�̥�� ��8����7�!�gѾF�]�&2�H�Z	"�tl���Ő�Pm�A�*٤����l���<k��a�Z,:�����{�4_�w/��b��C�+�QV�ρy5�{I����z7������%űt�㛣�y��Q2����3#, ����,�b�ڽH���� b
ՁM������]n��aP'E�.���u�<oW_��a*Gk�|7|�y�[����K/(�g#�qc���qn������G����-	)�dݥ�-�=|��[���>a!��U��D
����d�.�s�r�P��T(x��p�lA`��-G�7������'O:��M��m`�匉��<K� c�Dތj%��q��j+���n�"�P+0���C�*��)��Q14� �ng��]^_'M�֝#b\i��f�D�|��$�>+��d���wv ���O��ו�&k8�I����*�����C�8]۴短��ҷ�l�OC"�ەSsZ)rAS~�����<�!��M8��;2��� WXY_�nOHLEm��*�Ti�iD�>��L唢:g�Û^� ��,���8��$up{��#����$G�����@�n�:U�	���n<2���K��i�c2ߔ���c1^�K|�'˱�l�����%�cL�JM�H��@��zh��[L�}+�������B�Ͽo9�eV���q�˰gW���n=>�F���Ci-ʞ]�eW?i�/B����ñc�`0��=Ω)�ц����轏�-K�顸�~ M�a6~zt��bZ�� �ŨSQ1q1���{rt����������y6Y��+�0��L�5<.߱�<�x�M]7:K�0�z�"�'���rHj�����g`�EY1�Q�+>y|��_�����)ȕ��1�Xo	��t�.�X�����i����!��?�nN�U�>_�*�S`=��Ļ�Z=����z�v;H�)8�j���9M�rHÆ��#�xn�����$bǺ�a���n/¬�������c��T&�jzT�sUb\���>�\9%a���;H�?��7�l|��IY�8�����
����Ή�u�4P����93~��:��K��[fUO��pZ����C2��tI�G�B	����/##RЗ�}4}��M��r�;�X~��w5{��΄�x���j�P|[{���=�/�Å��~q��)�e�zy��j
`�{iq}Z��9��է>|e���Z�0f;5֕��܉�Ez�ڴ&H��cV)�s/-`�����$�����9U�#��<o��p;]WFw��]�m��_!Ԧ��"9����g�p#�������5mM��Y�x;]�M�-�I�n��Xh��ik���glLU�)k�r�K��ڸ�6���}+x�h����e����}����|�iKhve��k�`��R�v-EU�x4C��CJ$��=QJӟ��/�8��iO��6m���ݐ �eP΄��ڽ��\n��Ҙ�G���o���fV�vC���ϵ@ׂ����i��7�K�
-�@)�G<uHG	�Z���㛑[b<����\�����*�K��^+�*>at��x��^��~�h'��������͆M*ooNC_Y��WL�]�J�O�����E^g��z���`]���2��oBnq������?��#�G*3���WWewN�/��oV�o��>��3�� �{��S]�P�ɮ�=���{A
�j_��G��ϑA�~?o*�q5����e��Ƃ,������'��rg��/R�{����?~�p����Z5�go��$�k.�3b8�����l�*_�dL�w���Z��S�{;|rDHOO�I]>�7
P*��L�0�ETo#o�J�U����|��͎�������]���H9|��� �e�����s�x�1��Pٔ����5NC��U���qH"B����5��_��e�A?��;:�KZ����Eo�A@Zy���e*ͩE�e�tG,w��/����ǿ����Ԗ�8����/wD`����.�t�>�S�����)ٿ��{;��f�J�=B����;����(�G��?�%2� ����N�U(��t��sj�	q��<���*�|v�¦�.�.A�UUi��D�n��F������;l^�.QQ�A�]M_%� . �Ųm�x��I6֊,�Ј��� !�b.��l�F��3xmk�+���m�0�w�;��c�P�7�U��΍�zY�
���b]�>�����bI���G��e�`�~���.�t�ɪ��_Z���W7���@�R�2��XQ�z(j��bn���(�-_�wRn��_����&`0:4�<׫�N.�7��tq���f3V����V�;��qm/������d]��JO�Y3+�%�����߿=�C������~k��ģد��y�Y�ךs#�f	P"�e� �co�D����=;\��|�G��T 3sD��$ K7s��������4�-�(��\V�Go���		��N��_��{���^��	�x(������z��>(��g�Ih��aҚ�:��r�/ ��c/G���Νt�7��ޥ6���sɹ2��*�Fd���Z7���0o�b8������l���׮?EN���|y�E�4�]�.�I����;l�oR��'���������Ȁ�3x0m��r?|7H���A8�-�z���<Xc��k,,}=���Xψ�N��НEEW���SC��Am�R)���a��tf� ��`J va�V��l�\��#JFX�: ǷZc��(5���;��x'���P�������I��Y��`�"1j����d�'k����2"JG�ǣ���SW��N�J�G�J/����9S�SOH�� �Fe5T}yU�����vcn�;ݥg%�ﻖ+��[�Y4�Y�/��O�.I5�e��&,ZֆX�i��4w�?G^��\�H�6�&�~��F���t�0[��;���Kab�=��8�TT�8�rJ�D�P��c9ң� P��|���yUN�:�j���j��j16]�����f��i�Ҍ�S�W��v�S\����٭)6�ٌ�Ԕ��{�1i�'K����<&�K4ߢ^��\���3	ҩVoL���Qq�翞�֒d�xZ���,�F�Y����R����N��r���g2wi��o����[pifq��f'�`�(ԐͩƓ�`"8������Z�F�����z�x���)���(5f��3'&�I�c[0w���K���1��E@���a,@�X���Q�7��1��k����0�:L�
N����d���4�e���ǝ]d���s����F�|���c�����>8�WiҴ�CV�>��K;Q� ��#=�s6��W�VV^s��G����K5�v��T�v�>��f�Ϧ<GQjk 9��p�-i�<�$4�=�i={�\�,.�]��HߒI��ѧhhn(�|��| '�K��9��eBsxv=?���L 1��֑T�_x�+C�����El�H�?���c7$��ooi:���&u}=e���w�/`\s���Z�I�_VG���Q�T�H���@���+��wu{�!�e���s���Os=#�ô�z5�@�q���u�<e(���7+k�{�jA�b�c�,���G�{2=��d3B�0�b���q2��s���T�&����+vG�$7��ё��dK6f���Γ=�5��3�]�i��"�p ��'��f�}f��
��#���w�vb0};xOy�j�Գy_�>��.��O!b�f�>��k�X��7�?+J췧I� 3G.V��A�6j,)�\IQν���xBJ��s��I�.�M�@kh� e[�YK��K��z:G���izT��tG�:���^�Ӷe��~��<Y�������<�G�� '!�����m֚�W_�1�vc	�li�ˉ<:f����eZ��8�����-ݰ�p��"�ˠi�Ux�~�=��veĘ<K9�F��!�_�ց��1
�x��u���F
��Ն�q4فAh	}���'�0���x�_#���>@�=>��<X��0KT;�K�q�[pQT�.==�&;u�9���2t��F��M�Yd�BI.��Jc6��O��V��ٍ�L��`�tJ�>	���M�xUh��-$x���u�N�d�߬��-6����E�&k�����r�5�IC���l6{^7 �g��0��G����,Ԃc/T�m-�|�� 9(|���*�h��U�5���e����/AtH���D���nW�e j댗"����qw4���{A���f�3�髲ݑTu^�͙��jާK�+xu1k-v� �WJd��!�G��i��� ���m?�Xo���K$D���G�ue~������탔��
������S�@¸z��~��l�r�v,�_���D��X�kAC��j�^ֱ��K�mrb��a�C	?��=y�KAx	={�)�n]1�4�zX�}Ǧ����U��?$�h�����{�.�i5~���Sr�/F� )WA�b�H$��g�Ez?ʃ%�+ϣ��\E�^�iD��<���lvO�)$T] �%��d|��SҾ#�-��=�.�R������u�S���ݭ���$[e�b:��
��/a�_��fG�D;��vb�?|a,e�ZZ]�~R��C��!�ڬ	���0	�Q��78�����A�l�Z1<�-禪
T�I�����$��/�0X����w����@>�+ƛ�&_b��}�>L�1�;?�Y2Ҝ��)��GU�� /��5���H�e#(OR�������d^��p��7�0��Xe�D�,���'����:�^y
�]��.�2�ڪe�z�{�>�yz�����E�%y�a�>��!~��Q��$6:�~x��ERYb���`� h9UC�}O�֬�L=&�OX�_��ƽ����g}A�I;p.�.��V�������
4��3>ؽ�q��?�ҥ�|��ܬx_Lf
�)r&dux�-��Xh�s���|��}'����Ef��~F����hQv��j��Jx��3t#�y��4�F#�k?[J�p��	�#�D��I��T"�ѹ:���_�x������n���{�iʋ};d��|��~���R{�������0S��NU,áQc���&4;�1�������'U1ɫ�D���;#��<=�{���AG�w~�'W�������4l�<^�×�B�]\|7��X�陧E9ߜ%(ܬ�fk����{,!:�MI?���f9T�ƾooﾻH����e���O��������&�ţE� �Z=CZ,{]>�O��*U�+��e���U6ى�~T:�,�6�>
�ey�M�!W�!?~lp��-Kzh�L��^����N���!������f��]�ܑ�j,���{���8$�f)�s�Y"�������Q_�\=1�yS�ht�\�!H�}�N�H�2���Ӳ�<�n
+L����w�AuL��nz♌����2q@�*An$�s�Zoy>�I��4HT�Y);͎�� �~����2r��i�2X�hX��$~�|�޳x/p�h|���*�G\Z��k�<j�V9�,Z�ȷ}�BD�$C(/4Ƈ�b��R^έR����\��&����:[�4��^>���MZ�@��muM\�"1�h���I��^D�����H�6&�bW�1�@	gFQ��A�n��q�5��3��O�?\G���%[�^��5�C�_�TQ�٭*D����^K�t^#�p`�AZ�m�Z2#�p�sa���c���l�"�FoA���-?�Zn���@��}<;�jQ�(OF2�X�~���Om���������5�r����l)̔����U�R�鈳�I6��"6!��:��/.t~2�v����>��R�f��%I�',������v���W\!��;k �a��EԞ�|='���>9j�3�I9�������x2%����{3&!/�A�u~1Ӈ�A~�z�|2�,�����>&��4#����~LӰt��6_�L��XGV|���Sc����7���>�m�PK����gR��s�;�6�����A9ߔ- 1����1��)b�-R��0�\��a	���9�xH�����������1�05+��ӽ�������=US@�*s(~u�Z�WC�SWpe4�R���*��$�v5�zE}.�}s?8����bьj��;��;�~�f�~-t��o�EAV'xH��7�Ш�1~|�B�U��Tϱ[�}����;w��B�o�	Zf�\P�z~#��z��
k�@,`1).o3�t�O�����K%�t#B��߹��8~HFMUj��UtszOL��4S.�ݗr|J��=wbi�j/�%Z�����c����,�ĎH���i�x�<a����_[s�C�97�>7ܪo���T�B?�� ��i���P|�G6��G��m��P�3w�������v�|����v�wS�n�Ê�'�G%���rz,|��#5`���(�X7��{��{K}�/Ft�`T�x̝�KѼ��#�m���N�y�ѵ�_��x�c1�3��pL����P�M��OR��(t��9�|l��؅�N�<�^g�,2k��P��U�t���Mt8���,��cO�1���Ҷ��s���v�a��j�)�h5s�ɠ��m�z��-a@rErp�~���7/�Z �$���L[�wr����S{����2uT~��US�h��_��(q>
�~u �2N�.�s��Q�5�3�f���!+�#��T �����`5#Q!����b�@���g��5\j������|iY�Uy5VjX���ELR�V���#�L��p�P[�T?X$�D�G���?��/�J V0i�&�f�-`V��T/]z�3�����mm'RL�D��w����w6D�Ća\�ΛV�<��ٿ$��QĚ8��U8�,&Ch���h�� DNe;���Iɩ"e U ��\@���[|Y]��2-m�4�TŠ$2�.ԖJ�i��?��߮\��uCޡx����巖����}8�l���YF�T��t����*f ��Fp�GH�I�]�&�PL�M�י��D�f�X*����؍v�:�yP�K�U�����*��P�ٷ���xRW�ޟ��p��h�j�J�~8׳����a4���LZ�Bz������LK���C[#H1��5"�I+�����ˡ��	���R"RU��P��5)�/�oǋ�[�T˷�M���A��~�Dj����"����"��ŎU,����R79.�)�G��s�i�"�O�������#@�j.�O6��4Ʃ7D��%��)��L��h�U�|9�>��᳖\H�5����̘���57�T��t���f�NuE�rG���H�0^NP��ƥ2�� ��A��@�ñ��@d׮�(�R�7{Ǡ�n���x���S��H��Vb�iN+9�D�9�h޽���ܥ:�e]B`��S�5^�/�y��a�������[���d>��S9�"V�/:����}�)�<i�Q@c!b<�P'�j~Q�<k\��ц�lB�rwX�z��ܛ�<����d�.�
��e�ݡ�Ù����٨e'̶�`�
D-2�檛fB"%�&:��H���)�Q��v/��D~Ph�&��3wR�������M��~���7[
|?�_���;�?���n�)Bo}�A�!p��[�J@��̣������q�����E,^��ۋW�!��ք�v�F⑯�F�s��̛֤��ǟ7$���QW.`+������_�y+^WL�=:�Ա4%F�i>�걥X�	>>�G8F�Ɲ�隊Ap��d��N�/����fi����s�qJ���"��43�c3�� ߯A'"<x���E�?��^�/�,Y�/t?v�_ �/�sH�U�P����A�[����� ��9��8���*�+~�u��������7.}�	5\"?������g_f$2q�1J(�l�}X����\�Nj[}{�B˼�M	*1!%M�m��"bR�z�T�N0��MH������V��iM��:�W�*�� ��
H�(C�G̹و$�9n�c܊(b	:
E��N�
���;����s��k�C�+���S~��Ҟg`���c��U�xZ�!}��$�U��{�y�{��b�g�h��A�z;�n1����UJHx����C^�c�p�b4�ٓmI{\�7��5�W���h�q>�B�U�<�RL6�|o]����o�F�t�O�u2>yQ�Ɨ/`^�����IHx�%PZ>�;N����Ӕl�_΀F�4l�� J�-��LU��1�^$X�xB�:�T�l�J��kE��շ�)ې��;x����F�5���7�L��F���rT		��+Tm^U���j��i|:Y�fG�.�x�m`)QnN�d���d�
�mK❝�w�k�K��ư2�6zے�d�l��ԯ�_��˞a('�~��5|a����i� !v�-=k-Y*�l~�*��#�t#��"J�7Κة���S���xdĕW1b]��6b��Œ���E_։��׭��O�>u��\�����)Ҧ���;m�$����O
"��]�<&3�ldX �~�� �b�/�8�f�S���wյSA-AږU��D8*ߚ[F�޿N�@�'j����E����i(-��~�=�jE\���G�/�+�l�W#}��������P���]�*��9�f˜����_ �r����o6���m#/G�����n��/ O�T���%Ǝ�jf*�,��%�c��݋X���-��Eݎʎ��D���B�٧T��p81t�{%w�m����X#5�&kl���t:?�k!��"D��w!���h@ߺD6%P����m��M���?�;jD�e������7-�Dr�����\�ԙ��3�s���BDF�)H2��~�=#M����;*����t/�x1�4O>��7���O�D'L9��0-G�ך�Q��ȴO���:��q'��4���VCZ\t6*-M�Hߓ��\�8oN�h�����R�^�ɋ��3q�[I��2Z56�Y�@�����Mx�Vv���E���� )7}v׾[�kelt��jVy�B��h��F�P˲�i�l�.�P��gU:�p龵����O��P]��$WfC7�'�b<vw(�'i�^mU���eDC/�Qe���W"�S��2�#κ:�	 �"(�i|���O~���(�N�E�;�'q�<�5�i�W�8-g�Q��;�ǔaܐk,�!������L1������v���[w�/G�!�Yh��寉l��k�"�� g(UVA)YnC/O��|r��$��r~q3�~F�2u��%$ @�M���P�%1n��_�u�5���/KRgb���`� oz�-��4���	8�M�>�*���S�X�����I癉��p�x*����,�HiuKj��w�N^Ci���]�ٞ��?�ЕD,��E��AD�9�`V�zQ�3��u��A-���#R��	���!�$��6��uyn1��,�6�2^6WT�A��p�8s�ү}�Uʶ���2V��d������MP�w���x_�w����;a�J�PS"�ʾ��	Z�+Hw�D����=�X/D՞e�[ֽ�*�\��H�������ڨ>}���)Ɨ�[hLz�UN�:N~v8uGrzư����K���'����(��ʾ���~p/.*\�N�)�l�qVO�����2o�D��%Q�a��#Tͱ��Bé��Z��G�Ѭ`f���?O�J�r��]:�n�l&��<�	�Y��#-i>�[5�����x��t#�r��Z��wpE�p�'�:2�r��r|��{�񥕦��e�W���:w�y�^�7�O"����_DoL�2����f�=��d���w��o�vv7n�S��Yfy5`��有�FFF��y���~PK
"nShl��ٟ�[2��hZlY�j��B�[����w�ʿ��҉#�PQ����+�vd���S�kk���+�����[�s�L����̣�Ai��M�N��/.������}Ao U�lg���7`�y�".�vO�	�����+�M~|���\�uV�T�əD,O��%j^����Z(�%���j�*g���U�]7���������5mvǸx!7�ҧ�~QL�@2�@ʒ��)�/�OZ�0�9Jp�Ҭ��I����ʅ���B�ave����!"��d�̗
�㏯�:8�L�zztB�#׳�*i�%�)��Z��b
(_M3ς("�͸7�ͺ�%�ǆ��K��&����i��ᠾ�w`�-wBT����g��^*`5�8�,�9M��-de�U]XD�$��V��T��|7'I.<�#AP�K�BP�yާ_��\���f��KS�N��c��V���ޅQ\O���̠㧞~?�9:�ZZ�HԢQp�3�m�����"�����#��d���a]L�3��f�p�%IC~|(�~f��U����	�H���	!��u3sG�q'эD��+�:��ڡxG��`�/A�1�-��9�C����N���w.�����E�=!�����1z��W��)(�a�3����a?aa���V����7�k�������5��Yc[hQ�(V8B��*�|���b�����U�;]4O���'4A5�F���r
�RʳĜ���@�N� �����w��[��p�/�k�g#�A!71�p�2���vQ~p2��#ͪ0��f���Χ8�����Ǉ���𾂁p*䍡�iP'8���K'r/"[垺����6(�g�|]i���6��K��f�}T{{|>b�:r-��V��ٕ�7Y��]�z8�_%z%��D��K.~ƞT�뇯"M��}�Y�r��rύ/π�b�������MN����3 E�-�=|��4�)f":>��ؾ�$��`�!�"f�U-�ح�=�s���+ߛ7���>MZ�<���кC��Lf������?�����s�LI� "�.:��d���8�{�5�4�\Hmh���6���D��OT��i.��������Yo���J�>cdd�sԻ�`����]
�Mo�A[��3++��O}�b,tb�v=���nL��x�e{�m�_\K&<�@+���\�,L���X����ғK�$h�Ql��F��� ?����)+kK
֙�`�I��U��Z� ��������,2h1����Q���ʉ�	>�SE�E2e{�!]�Xɐm����f��L:C-� ���P�S�)�O�KAqN@Ul�<��H
3� >��.������]C��œ�I��s^�'�=<a>���L2���Z�h���	����|!��P�p�1[$�Z6cԧ
ԧ<4Oͼ^N���wKy:/`q�ݱGgS�$S��5����祐�q��I���7�h�q���9k�QI�E�$�B��j+��=���s����[�K߾����7�(PbY�#7uw�^�j_�|�x|e5��b�T��d�J���Mc�<}��ҝ�%j
�]�+�|&;/J��h
���;;�c%Ѐ!v��!P���Uk2D��@�f�K��:�F��>���md�`q(��d�'#��7k��o�w:�ƽ�v]a�Ӻ��uԗ�J&��N�T��<S#��ud�/��2���6�;��Պ��&�s�H"�A��|���I�Z��x�M,�	�H˓��N<��+�KW��S��x�?^<�u_"�/�zc鋹zK7Lwm�����%!Qf���e�R��
��uyI�4�kn�G~�X��;(��X������V��\N�u�h78�=��C�wn��(mre��߯ЌXo���B�/TsM�i���Ws�>�'�{�dYI���f9yj��%Rd��vb��ԇ��k�����) �1��CϾ���RbW����7Ծב�N�W�o��ٓkLSa�͒3�$�@kh��^P�tG�����Ɯ���2�"�h�m�\dm�h���T$���������y��cE��W��j��P��sv]�U���&^��b�S�#�x��5t�� z��J۱�v�d��q�Ҧ�[�Դ�n3�n87}J�О
��?Y<"ĵ���;�Ew�|��6�	1��j;��~�ֻ�ĕ>������ؿ|�Ŏ��5�n��=���#<7��E�\�%�y>�tv⮬coU8�����M�$���|�Ϲ�	�p�'�
����ҝۘ���"P����9������R�!�O��D��l�1�u�ݢV��8&[322�bV^P��5y�=(�����k=V�t��*�W�\n6�Mtq��jf7�H
.�r!�{Ս1~��=�X�	kX��=SP���Y�S8~>Ŏ�Р�]>T�*�{aɠe�A�?J�H��h���j\�������wh�o���WG�q���1$2>N���|���&d� l���厺�<=Ki�ewЛ'�M�N���zڝ�HF��{�˃e������1���c!�ڋ��iIJ�鲲���|#�޹����ţ��?��b����)�kò6��v����j;��}9�c�+��g���I}���*�6�U���z�̱ߎ�qf���)�d9�	��	`6�̿jK�X�K�0Չ3K��#H^�����{,O]�5E�� ��u�P#'1ٚ��x�42�q#�!��#�&��|3��YJ=�v!q̓��H�u{t��5�dm�i|cKr24X�7F���vϻ�nS,+�$�P�_���n6<#R�����Q:��\L�#��c"�NS���O��޶�}���HZkO�/���h���N��d֗_b���~���ON�@Hw�+���Q�+i�����	����0���J����i��΋�j�;�Nr/����"/h����x�~Lh5��j�Y�<�ک�f�ܝ�hXO��K����Yr�j���'N�s�������f���Gk����)��9�� ct��9���{��;����~�jӢ]�؜~�Vcp�������(��� �l	�O;98�{^���sv�9�n�G9��h[Q�"�Ԝ��I}\�x�B�F$��[��+�m6��g��4�=r�&0�|��S,+_V%�c�.+�K3zA�X@�����|����T	#&@(�ⱉ�0�ʙK��DB�7��%����"�ZP�ws�����zDAT�ژ����G��d g�=V|io7xH:��3r�$s��zn�%Z�
4<��x�"�~���g�����=��'�_��CT���(�zK�hS��d����r��+��6������뺹����Bh_(v��L҅#W�5����!�1�j��H˦+@鴀�������P㳝X��x��T�(u�93W�3����J�0#75��v�)b�Ty)SR�+�lC���b��>u瓿�D�ւ��B�\�}ꀁF�G0�Mi����ީ���+��=c���?P��V�Ua�V�]Z=��7n�����O<iqz�W���y��(}��	9�UCh��0��p�L]���,Hi�Zʥn҅��c��N�إ�0�����(�u��M�Z/�K��k�� �����Z60E&�i Aٛb��q��j���EJ	�*x�T����LF�^P�E�D�i
u��2������ 3W�$0 $�g���2�l6O��s����˄QcH��i�B�����T{��x�� 4�j��+�Y����<�"Gy;�1w��HG*v��p���Oxw��&m����P�F�	{����ݳe�ڋ{0�BW#���4��D�M��?���;���Ms��"�v���u��[�]_�S�$l*l�M%R$��mrL�(�l2�&���^\'�x����\�� -Up������X��M�bQ�\	T1���������J�A(�!�Ϙyl�<��sC�?�r���3)��5�����i�Qc+\s��P��p���(��"��{._�U�8���(���s� Nì�x���%�Z`L��A��F��X�{^����Z��b������y2�/{�kc+��w���O=�[��K�ĪK|w�u�,h��j�Wa;c�J��8M��>ݟyxL�Ym1V�{���9%�7I;����P�J����^�s�0{�_�a�K�d��*N �	�j�**�7L �^��tKz����R��L?q�R�������ϟˡ?�f)AN��ab����"�d���w"����Z<�`8��ES��/�*�m_`7yI\K���L�A�D '�[=6���w�7�;N���S��bccã�w �fS�W�6e�Bqp�%5����?N���8\��1oY�j�,����_U�ﲿnm	��~9]=��;�fң�������zAN-�)�3B?'�m���x0'������zJ���#�|�%{��v���� m%�MǕ�J��G���&�6Uj�&vi�O~~`�ľ��3����P R�<w(�萋SǄ� �jZ9ׄ����@7++��1����bT����f���x�P��޳ECcS{KKm��5�
�7E�*��b�EC�Z��b�Hm*�����=��s�'���z��x���R纰�K�u���9G���ڸJ�"���$W�m
��D����F>��ۺ�J��%)LU�<�nn��t۳f*�5������5wP+v' �!B!1A�:�Ͽ�'��W���tf��b&���J@�مnaXQ.H�3�J�gCZ[�M�x�� ��GoC�����[5������?D�3Y���Z݁2�-�L-?�x>k�ϷRR�lv�y+�
���X6�n��c�@9���h�ggfTe)��v��H>f�k{q���5����$9���ɘ�&5��zfq<�����G��z�-��A�����;~�Ek\p��hߪ��CX�{�����8>�c�Ev�<�&0�nx5W����1�R�ZR�G7�������I*�`���Gʖ)�9���q�~W��w+�Q����/�������aI>��n�m4�ޘ��HFM9))ťe�G�p�����dsv6���C�w���̻(t9(��υ܁��P��:{A-z��������(��nPZ�f`R��3������K�{���WE��S�6�|O�>�L����������0��i}�8�c���~Js��r}��w�X���/4]U���p=#�GU���9��R.j�޾���ҿ��N����zP׉�R��0��{�,Q./߃�c0���,������r��kЖ��H��o��TDv-�k�)�<�T���٣�&��4s�_j��c�5�B�������K��Vu~�	�7�y���B0]��q9��\`��V�<���Lu&��R>����G)*,=�C���:�d
�4b84��S��UN�o��y�I�)1&��aS��I�U�r@�^�/Ԃ�D��C���{�xu�y��[�ąy�%\�P5��	���k�-8�\|LX�E�q��� �{w��o��&�t�<?��������W��myq#/�a(4�T��j�q�バ��l�OL&�H8[׃״H�80��nq�U}Q��r���.�J�?�&������k�����J��yT�Q'v�oKӈ��rh��4x�P,�3:����y��h̚�q��Q�	$���}}ҷ�^��¦�[C.�n�tN��̬L�P���O����'ڲB4fL;f�ķf<��C�<-c�N�kl_I��~��8cx���(Ó���bl˫��y�@�h��Z��=4�gxg���W���m&�$y��;�DֲҮ�Y�ղ�J���6�_�3���� %�0�.�����t {��˿���@K3F��ucj���z[c���ɿĞ ǾX��	��7�[�h�W�RAeON}hXU�3�:R����`�ɸ���.��J��R�S!��ɐ��UǨ��BS[
���l��nW*�P,k,`�j���td��^X�F ޚ�HFe��0��7�C�阙S�jJ������<
�g���l�������z�x�Ŝ�a��+e�N}�0Չ$�IM� �4k��*��CD�Q�SGr��ʟ�zZ���	f��$?l�܏�Ԃ>�ٰ�ڳm�����G�j���`�syOOO��֕u���ӭǀ�����?
���j�S��e�'}ɬ`���~,\?0�����63��<wh��
�?R���딂dhLx3i.�����q�4�?��R�(d�ZBL`R�Z���Ҩ�و�1��� 3�7M�v�:E�H�u����p�Kŏ���v���0%9cĖ�0 � �Ұ��УD;{t�! � �D��N9KL�������AgUƱR&�K�"��؜*�[��-�7���+��I9�f2?�U�7���~�_�z���u <��.���N�?>F�v���T�e�~1w(=d-���UΥ* T��lbY,�ܙ�xQ9���7t�ᆎq�t��<����,[j��L�W�S���h�u��� �� oU	�$r�nFah꓅��`���F�����N��H�^���ά��c]����.o����{F�J_��/Zg�W]���  �(W��C�����{��z��=enu��j��Bџ�����F��i#���X]�x;�FX��m�kl$��鐞����8{�!��z�O��(�d�?�		�W�2�孷43K��z��qx�FwnQ�oHG�D�rX�8YVɖ��:B;�m*e���f3cnZ��I���0� q��q�XWu/�B�u�)n����9�Q�ft*���A@&���������j���1!�]N��-e"YHk_:��ٶ'qeZP�?��}��a�=	I�
M鹢c��n�:�1PC���Ӳ,�e�6M��I��p�(^JJe��x�|�o��T��� Ά�H�J��E|jBj��>����k��:?�o�i�*�i2�{���e�d�[��(�P8pf75$�Hm��n'u�a������j�C�h���V��q�L(e�^p�����p�2F	.�X�k=ٌ����+t��_����/�(��p�h�"��ǥ3F4�:��%��Yܧ�
��%S8!^�&�2�ޞٗ�b�0)��Uf�jH�d4�l�t$yc���g�0�qRz��8�rCa�M(�������S��dwW��-�(��bba�x<�$�d��FJ��Ȼ^�~O��%ѼTvL�~�C;�΅�{�w h�wޓ%3�s?j9���6�46&\T��WJ�=*�����G�t�4Y��o~LF�n��C�r���w2����k�*�~�F�/��k���J�ꯤ>��T1q:;:��v���y���L^��s�U��FP'i��X������f�y]`͊$�;�xw�>{�!�W2����������[A|}F�+�ݨ��S�)+Zb�| `Q�7�&b|0oր����PM�囨�IW�?��H�_k�	�k�����Z:�$�-T��w����5�ސ~`����QN�D�GMN�����6i��<᫁�ݢ��[#'����FT4X��=�|_[������􌍘mXN�;㘄F�Z�_���j���茅��c������2�-}�)��T�~�8]����߿�"�q[�J!��j���L��_�����2���>�ٟ� C��y9�.�W���sV��,���h��fU���9�vh>}!���Tκ=�b&64��p�efI��- ���	������$֛��~�\�����r�(5���c�h����	�px��s�}��/g���=�e%q�݇"�Ʈ��qD�B��7$%��󧤞f0�B�O�,z'���kIxhw�����ń\7�yj��1Slņ쭨Zrx��`��xefF�2Td=6Yº㺰�O��'�����o�_��A}^P��>�:��+�S�A���r�S���896���r	6�;ODSp����9���K�!�c���!�b�3���\���./9Yiڱ����~�=�6��O�#N%/��M�������o�֨��&/e�9^���I�{����E*(�LIjh*K7�̠"s��"�@Ս9�>����BY�)��# !ߛo����P]~� �����],8�NX1N�Fk'��/��]��D�٨��N�02cLN�{�[}s����Ab*��P�����:��{�sT����w@+0���K�������W�W_��ә���8�(��׃���/��O�tQ���m(�T �$�L���Bu����<�/�J�
�F�O|�m힏�����6�F�,{�^$��e��C��q�bC�
+�'�A33��i�'�: ���%nli�x�n��<��Nh�����w
�'}��n��;)�ڔL�P�-��u�|9�$cџYȦ�%��0J۞��DL�$�����(�5S�J4j��!�n&0g��f��R�i�w�:��! y˓q��l��r@B�OZb�dg��5W�-��]�p��7yfH�lz/�)�ZY!�m�AU�Ő�)Nu��2��^?�OJe�������/ /���7�Dg�:n���Wà�$L6�����ԙوE*�܂\� �1 �s�.P���򪰮\�pC�N*�1:�u���$��7lrW�G���M�[>�%��prk��C���Z��qw�KlhH�هO��;��?YJ1pp�t�wOi�T5e�:{��"�Oq{�Y��*e��!���蠿s3�@��ZK����=��|��ZeA���#F����3� o��[�	�~1��	+����e&�w ���:dI�?��٪�^x��KRi�g�����TZ�"_\q`�')�2{o����bTRD���aA:��ؼ���4�у3?c(�,
Z��
Oxƻ�a�ơ���d*�'>IS���o��
���?��,�W�K��-���Ů2M�l�&?����>�KL��L��5g�,)|�~�bLw��U���27���XV�ys��Z �تfn�K!Y�a(�����dH���l`�4�1}ۯr���s�%O�S���^W(U5a��1ܡ��.=FU�������(3�;��p�/e]�1���B)�M/9�V[��\ͤdm��t�*��-��K��}��m�?��=���(�yVD�O���O����,�;�~�q����ך�֡y	M�2]ތ�;~T����=�|��}znb�5,7�J]&"'���	cY<?g�����b�n?wrzZ���~��Riw��E��o����:H`�k��(M����?��k��,���v[H�P�G*�9�wd�ށ���l�Gg���G��-�%���E�;�N�y_>�,TXT�D�v�5�$�4��7��ʹ���G�TfVJ�Ⱥ:{�����|@�N��1��>q��V!� ���ZW��ۺOJ���h�!E#�x�ByM�x�&��ݞ0$�DZ�D�|��l�.�e���B��H|=�D%֡<�<P�A� ��|��&j�h�Z�FB(�7�/��M�E�є���8�e������$ֵ������%!2�+��}hi�fg�*R}ѧ�6�~�o���)�{/ɣi"򥇛�� I(��WV:݂�a����0���R)4X/�~T�K90��3O2��y���S:��ޑ�C_�xMF4�R�00�Fs�K�F�e�E�����G���0|y�P>����=Ψ�!�1'��­+�+09L�^���R��V�����]<;X-e%_;��+��<ͬ����$��T��cH&�q=<|7R�c���((�d{g{Ն�/���}�l<R���IU�S+�c(���<���er��7��$v��|�f�v�;�A逈�5��p��ݔ���gޙו���4�L��cg�etӳo>��^C���c�+>�o�����4���XNQ�L�%DC2�Ѫ�;�P�>{3���΢����~S����F�x���$�»S'����!V����նm�f�oΗE�je*t�<�|�8@�9����&���dr�zQ�Z�rdTe�Ҩ*'��U>͒�8>}ԓ��/By7��}@ݘ�4���ap7�y��ޑ��j���U��Y�03ÿn�I�-���(]�59��X�A�@?�{�+8��-��!�0$��%I���rCa� ӱ��s��������:��Eo�����S�,�h��ς�=����.]�7"��G��V���λ?��(���0E&���Lx�O@���}�-$qʝ��fwX�[�E���t�V���U�=K8&%/#h��ٛ�L
�}ݔ�w�|�o7�d_ɭxV��;Q���� D�O~=���)��Wp@�j-Od�[�
�H&yUWW�i:[�*Tq�#��"6Haq�m��)�s�58N�ׯ����=~��p:�"v҄�n��8W+���H��ܯX9���/X�>c��|2�h��`&E�����#F�౾�]�i(�~G�'l����R����K|@{bxA<z>��2�N/�����P�bp4k5L�{��Q��~+g^���-��M�y��B�N��um��C��+bZ��j�o���(��Ϩl/�#����c�^�[y9���EI��(���찴��FNY����"�y��T���@:t�;(;'2Tc��7�d_q]�|��}�w�_T'����� o�'~.WTF`;�9=?r�50c���ꜹ�=A�ІYGGgr�ƅ�V�������ƍ����L�^�\��"٧[���D�T*[���1�K�y�i_H��>[���ǝ�L�0	Gⁿ�I­?^�*Sη���܏�?�O&����_c�_�� Q��.b��ѧ_i��26��3O>�,_,�rl�{��T�IІ,����RG�c�i�"uSf�ۈ���� @�A������k��u��o�'�~����=��X��*�3Hb��D�sL?-qE��j��+}i������
%��w&���}������'�^�og�2�>��'�Z.�W������@�k��L��t�
Z��}����
�������D��V���`N�^��|"������[$b�e\Y~O�^[s���a���Ǳ/�W��-��4�������i$�_o���|�`����������u{���ڵ���*��;�{kKt��#����7�W���e6���r��2Z�����n�57������ß-�eK+HҀ!<CwNC��B�w/J6���2��>+��A-ȱQ{����c�S��di�/�c���yT��ߓ�'9��gAo����x*��r��v�꣸��u{�5a}g3�ۦ��w[v��֬r׸J�
�z�d|I��D����f;q�ӟ�$�p�=6�'�b,o⋠ٺ"��g��5b>�HΙԭb#u���ɼ��T
]�����}c���4� ���U�Z̺y&}bH���"
��2���%�m�:�����~nzx�ٻ$y|AdE8���-��V\���<��pT�P������	�?��JQ�B�|A�U4����/��Y�H���.�yE�%���q��뗛��<�0������]`�O�������s�"�1j��؈������V�ݚOt�����/���G���P�y��-�k�H{>&��z��1cLxY��@�0��rɐ������43Sw�7��M#j�ɽE�T����]VN�������5���K��#ҥ�͜IvVLJ�&Tj5��$C*)QqG��<c4�]z?{Ӷ�X�B�U��V�I��M|�0u$w���}͹/t'�kV �k���	�����W�Woh�D
��0�F�'P���PLq�+���'{��=�i�N{k:���
ǈ��Tu5y�(o�����ns
��2��n�_m7��{ݴ��-,\�D�O��Mlj7���9ڃ��9Ed"�=���(	�Xy#�G��_���[U�5�;#^c[zL����RW�@�y�Gq=s�$C�,Z���X����� ����$����(c**�� N:��a�7��qhο�6��Y�Xfj�R�Puߟs����£~�E�3�Ehd��4n:X%+=?1Rqc�J�ņ��e�(����a�%Ki 8�a.=H�"NJIsc����~Uh�:����#�\� ��Ux�xN	]b-®�4��L�MY��V� y�'��Xl����Wm ʫt��p+�\_�ŷIJ���w�L?Bm�#��,
��h��[h�5���I񝪣p�ΎM�[�uf+3��]��|v�ϯ�A�TK6�)��|�l��z����;�*��\�[�5����֦�IO�n��(��h�<-��rR�6O��(S����l:�Ǫ-��	�w�T�+�溶�8��&���P�x���bn�N)�zȀ��z0�1�9��A�~L�����i����z;�pܜ{�e�[_�p�@�Wny�IK%��8����mq������׺�qp	O�,�BL��|6��Ҿ����S�/��v�H"��\�%�f�-1����薂T�,e�� �c	Ty�L�N7�N�I�K<�;3wK5�W�v�y;go���|j �BҐB�䐡x�`�G�C�-�gt� ��e?�}:Ngf�=��Le�;�͉X$��ţ�fN��~��5�$Z^�*��j���)s�Z��<�jRqqD�yA:����s�!i�����.�X+�;ۣ]G"Z�������o^�"'0�wM�4�n��ax��l��<�'0-�*���V�SV��l���F��5B<k�n��di���/4q��C۬�_�;k�K�W�SuͣT�]�ܜ>h,�K|��O�Ǎ�c��d��<�w��X������
�����ŐǪ����o#�=Ľ�x)��^�٭Ҝ�3��T�����I��!��=���yj\xrr�"$�h�����*KX�)�x�S���D��i��|�'S��rpDE�^��"+|,�Ƌ-���`%.{0��μ%�ׅD��^���L�W�55Q�� �a��_k
Mma�on_c���z"�S".Tw� 끿�Yc��5���:<�Z�oG�᷸M�ieU���ԛgQB�TA`Dl7�>�KK"��l�O42�0��{@�bsq�.��ͅr�._غiʞû������I�f;h�0qC_��b��/x���o)�c��)��U�
	��9ŖbYE,���.`�,��h��)V���q7�8���1�$p�=K��K?0嬛@9�2��&�h�1��O6&��pj�9[�?����9)E�DL����$��W��LV�*�5��se�9'�C#r�W�[���<3%"��tQ�5��qKr^��p(]v�I��@�S�1b�3	D1�#+��Ա�%�+o��+��e<$.��6L'�; 4��W��7��/���u��L�~�5t�}�t\�>��E�+q--nr��q;�U�\���>��vYv�b�k�$��<Q����'�4ʯ� �[��]���%�D��O��\�uG9;���1mƌ�۞�`x�d�C����"7�}�'��~��3��^d9��;.D56����*�������ܫ,�A�<�R-�� 5�w[�X�S�8�r'˄�1+?Pe��m �;� �)H��;J��訍F,�gȇc�	x	�T���Ej.l�A�`J�c@mί�ҩ���N�1�B!�L�4�!�	p�sK�BK��tt��zPu��y�so�܈N:�{m(l�1�x	�S�t4������K�bɡ&�Bm-M���)*Ga)��iT΁�%n[Ԣ��-��oҐq�9�|u�����;˟{�*%H�z�%��>2�J����Nu?|�4�,��}9�eJ��H5		T��몷F���awf@����̶֦N�A;V�0P�������U����NߵӲ��nr�8�۽�Wm=N͘_5i�.���|��ꖹ��8N�x>y̶� �]2-��h$rx�q' ����@�>T���%�##�w��L�{��#��]/ѣz��1�r�DaP�F����+ܣ�c�W�=��г�s�=�\>�[�t��mk�:�i��H�yCO�t�Z��;N�^�r�B
�IK?�đ���_x8 c�|�D��{?�bP�����̩�:�M\��Z!�{7�H�R���5�w+/�!���^AAq��m0;+!�?f1(�T��튎j��4Z�<�N���+�8h�?b�F�l|��K^+f��F�Ԋ5���;5)Ì5�t-�{K��i����h��7W���sqtokQ)��G��O������2�rQ}C�1�f���h"�^#M�ՆN�$i_~?����>���3�Z��٦��ܜy���yR���I�TM&��k3h5~o���[�a�_POL�b�c�(ɼT�7ES��zN��fʓV��z��.0-F2�h���D���j��Y�z�~e�O��#Q�1ֱ�I�:�9��^�rI�_�Ps�97�י=e�|�]�%�+y	�����b�.�{e�$�8�ń]���SD��D�fq���l��/Rv�{A�KXr��wPНQ֕-�QH���u!���8	�_ڕ�`1�����O.�ݑ�^47`O�D��Q�F���C'�E�^�m�i���`?2�����ONJ��t�o�<��s���*&�"�yjM2�D�P�&��km�[��df�P3�E��W@�2�c�Ir�7k�����N2;��L7�m���_���^��ɚm5��^�#��Y��h����U9|P��Gd��q�~�F�yg�����JQ�@��Uˌ����-�uf<�{��ǹW��_��7�
�a,�cT��	x���U�k����-K
�D]��"��:���Y�-�.���|_�U!�
ŷ.�� 6v��.OBh�����2v��Ir�&�%�A�-8�<Փp��QR�	�J۫�����pND\s������)ro���g"�J4�p��m�W�إ��%a�v�	���;�}�͹�QEV3��C��,�"�1QJ���?~�0���-��޵����-x�P�5
o��Y�-��x0j�ن`WUG��K>��1/�K��8J�+�(�)�ЩHH���M���i?�zV�E��OG�<��W���E'���M�ڶ�&57+N���qA1p�W2����r�C�K�m�Q2B0ᝡ{�����Q�O�޷��'�C�חE�=3~%ڹ���GJ���%C���*-�c��7�n�:<� 7΀�j��Jr��#Ί8}u�{1�i�/-�v�ϸR���:$���G��촟1Y��E�廊DT��m�:٬�1\�6�/�=�a�A���+�Pj�-�i:�Q�q�ӽ>&7����gh�(��K��s�D���޳�F���s'i�~�fT"�.���@���B��z�hk(�k���H�hTꀼ��Uis::���"�H1h��1�;��2��`q��Bo������F���զ�:f٪��CS�.P��%�&��S��W�.b��FY�(I\ ��3��D�����Ricx�\5�R����d#U͘]ؒv�eď��5�#��e���.9��!����X�4�j���;��g���(�� &�����e�����ǈ��x�Zk�䤚�=��*�C��r<�Mb:GHl^����=J{(YuzA��Y`w�QQl�պ�{�u��b*vq䅛0|��T� sY�����X> g�q�b��DH��#���^=$A^�TJ�W��}1t�F�K|�j�[�ti�r���6(v�A �s�����tr�<�O��-V@@�t��`��XV�V�B���bW&�d�U��:'��n��#���s<��%�8�
99�[J�xM��îSn���x�<y��[�.��s�L�Nwu�q�"�8_Ν m����ɻҦ��%h�������HbE��8|�����꽐����ܔ�133�N)ۇ]�3e6!/ըC�����l�ݾ���_��/8��5�F��@��fb7�1��j�JF6]b���T��z��N$u�AG���]�1���H��9�T����0�F�V���}nyy�t����w89E�~��h�Ȟ���N�>�c�г�{ ����͜�Q�ÞRE�vg�2�����λ��퀚Y����'���v������}yq��b�(c"�f[��A�n�CJ~}�E�#G���	�>k��л��u�_{��6xt
����(t���\��P�y'ߌP���Um� ���爺@�٤�	B����&Ҧ6������Ц�(��.��y��ܚ�Q9N��_N\0d|��T�����3��p^bJH�M��9�j5��N�\�����͵��Vi�-����*��o��0����A�TTh�|�O�����6}֙$P�a�j�&K�T����c����DS�J]k�4B$ &N_U��	�^����"�(3h�+Ŋꚵ9�����X���׃�Way\#����<�@� t��օx���J�>B���Wٸ�V�͌�x(�����[AF�^���3I�.��}l%��s�hr��.j�t��b�����a�DV� ��ÿ�>���⹔eDhf�\�(�ȃ��Ke�$�G�9��x����M�����X����E�MI�QT �_���(�ÿP��=�{��Vug�X*۰Nʗ���D�m̛z�-��C︖�������.���tC1#͢�k��pǅ ��?Y0P�0���3i�Q�����4���%��D�j:<\�s9��E{�W�=褰��ш����ׂ\p�!O:ſ��E���>Y3�BPF�������ZόƆ?�0��vS�mmXy3�������f����K�~H(�>oLt��@��y�Q�6Y@��*Q�~�Z�.�B��:�l����Q�m���.�N]N�\:A�A�v��ob.��AX*N��D��ʣ(-����H>u��`�G-�3�a�;�xy3�i���͒D׿ ��K��o�y��M�T��] Ლ%��� +ٗf/>r\��h��%H�z���=�=��&���=��̳;7���,[^ ��Bj=r�����]���ɺ��0['�[������Z���]pRzO�{IL�_��D	�r�� 6"�#}���?o{�����*&*&5��8v�]�/�t_"f��K�R�v~��zy5���"����:��η�?�@E9E���]����b45������s�E�����<[l8."������i����@�U'��]/��#/��Bq���*����K��f]F�@��dknY��w���2�O?i�>1�x�~�����=e�T�1uy��]�04��⸤7���3�����������,���X�煛J�GS��	Y�:F �4Z}���G �t����������_���~�&����ࣺ��Ѓ:�0��F�H�	Ζ [I�2�	�Wj����(�����:����C{�u�P�vuEٳ��%�����|C�7m��:
^��v��Q�̕ʑ�)����GNI  /%�����s��?�A��w�n�=ĆB,�:��o���ޕ�������68�t�v�Gb �؅��?�=x�c�|ZL�����ҥ�/Z{T��C���ID�k�~�EM-e,l��?R�F�5U#r���4���c�ΌhE钀�>
�]M"@y��D�3��Gvl����j�g�V���D��R�.3n�n��
8*i��ԓ/��Zg��<Y�,��8��w�:�
��X���D���*}���%����H��(xB��A ��1�D���x\�cx���t��Ǘ)Z3�{�q�O���c?�����LFU����d��< �CO�%�8�j��/t�G�����vPP3�����aQI�qs�-�sPrؐ( �"�b�P��6:I>���L#i�YL�f��V9�7,��e���Fc���*pG��ѭG	�������{�����J������*9�u'`#��WO���'���ͬh|�yF� �'�<�̤c�����x�Y������_RJNI�e.�k���^�a pM%@Id6�C#�%�Όug+Y���(�4��E ���붾 ꝥn��}p�E�����%&O��	��O�;��vrPٰ�i��Y��f@`�����FY��XN�Q�rh�J��Ь{fy�	���;�u�M3ɞ���]M�(Xu�^5����*]�]�L�}�WA�n׆;�H��ب�-6�W�|��b�QiH'͢o����W:r[J �u�1m���g��-�o�Y'�@���	��[��^��3�c�~*W�k��\��S���!Q�gM �(���T ��OCm¬����*���7��_d,ٟ�d�k*�%m�D��@��$)�$Q�X�Mm�9bg�aa�A+�V�Ա7��h��M�'���6���}_.��?����V��)Cd̟��qW�t:"PB
 B6��5�'ǽ��d˔���R��N@NCuMڗ�В!�ј�:��81�R�X_��r��Z�ɘ2q�+b�!���?�OLiK�.��Ю���2�V�\KsfզW�(�U�\Şs�q�fn �G�xX����a���ɇ�KPj�������a��AH�����o���?��1)���:F�#/�؞�wX#I�����ep��á#w�q�eA��FiL����lن=���Rf����[��W��)K�K�X=U��9�8m�)�I�>IYg��������ǧ�����M��'vei���ӡ�����qb6㢒Z�i�9F�2^o�)��h�����{�s_)�
�����
�*'N�娵W�)jh?P��Գ���"/���AG՟�Օ�ˆ�1/M=/d�wIy�veA\�v��l{�'$i}m��F�wW�'�/SkgU�.�_}��q	 4��u���`O�g�H�]��Y+��q��a ��\ǚ���ܼE�������)�ȧș0�N˾lp:a^�!I��&lsV2���q�"X*��Jr��̾'u��-�"a���f�6� �=v�&�Vߡ[rb����J	�Mw��h�Ce����SqH��X���@�ܪ���P�.ApXX��	���V��34�c+C.���K��s6�N�擜�-��kTo������Iq�w�1���s�ċ��U��h�1C�=T����/���ǁ^�gr�]�cUZ�_i��6����ݦ�5N���]Ԅ�p!�Wrz��7�⟍vE4��NN&=Xb�u�C��!�~uZ�V�~'Q�*��f;�1�]�_�s�3�g+=z�z��f�qƃC����d&�4�d�@�b�Mȧ��Z(tn��7Ĩ��Xy�c���ot���>�u� mO�S%7�.�;/�u9�����\�Y��f�O��w�x���y|ʃ!IR�� S��D���j�	���q\�ӎ��ԏǶDuS�:���SS����5�{�^_�z�q��ݱ�Z��h�\,Q��9����?&S��F=sQ�z�/	~�"l��9e��te��������|�<�a[����¸��Y"���{�Q��ڬ�LUrh�)��L�;OS��Ν��м�Sk$Ө;�ۭeM�Q��"�z�&
ݮ�� 8d�J�@��Rn�B�<��ђd��͗�]�h���b%�'�b�C(<��Md��ɖ��KDu2TI�t5 X�SW�ב�|E��IR(�Qd
r�C&��b鎬��F�h�0Zb���i����5(�x��y��s�UX���t�q~��@-���[�dL����?~u=4yK�۶S����V,%��?YKX4�SBF�θ{���x{y���Ή���*���L-nlj�][#/Q�e�{�i�2�&�x���L���>'U�g�Y6�?���r+�``6QO���<���$~�HCE�ф7�8�O���5u\�~I��ɳ��Q����4,g�i;�b��H�>*PN���u-��0{F����͔A�P��=���|�+<*�$��_`]�m���o�y���{_�թI���iGHk?8�? ��Ъ�:������"���S�(�
=!\C�r�KiHꝎ�NI��$x�8�� ��Z��U)���B[�N��s1UBZi�%�!1pc>b�x)O��wg��)y�⮸2];OB,3c.S�}6�ؼ�Ԛ�]��<%?
�s0�$�����0�VZwa�����\y}�d2N��.�+o�(�~`���&MT?7�
_Z�|wܨto`���q�����;워.Osb��N��UVrf���~"�>�@n"�?c�����^�N����;�}ѯ7*��2ſssg4�Z��bQ2�[��&4a�s�7t�����%ԂS+�'����$|[���b�޹�uX��PD0狺���v� �(�\pc��y�V<3���(R�֏N([P5���a���G�Q�\�Z��Z�z��=���@9-�W��z���U �̸�uc��1xa�l8�Y>'o����Lj�F�,Ū1AՃ�@���v��-�E�W+�eX��A��fB��T7]2�X�P���Bq@Z�b%|ͱ\3�n�r��p���ZC�~˻C��.��^w�.Ŷ�d>Xܛ��H MQ�ot������*�L��z�&۰7{Љ�c�3�K=aqd�o��h��h(���E4�?�+�z��.��*zsQ=�v��FoYmqz�r%?"�E�V��������Ot)�|����c�����X�{[ ��ښO��:��Y��޹�I���]������2�q�*u}�}�����պjws�;���S�������ꔼ������we���C�j#�h����p��� ]VVʛ�/{�(�S��.0���L'��P��'�Nw�7g��V�ؐ9�e��ǧ�6�gęwC�uFYQը��=Aw\�Ϸn,͡'���J��oB�{^�\��˕�ׂ�QQ�/Jji�o߳p=�����`^�Mj(l����Cmx�d���;v�����|I�D8�1�ZZN���𫖲m��u����5i�$�%��B�%8��5Q;��6Z���k>�.@IQ1
6"��"ˮyw�sy�2|%�߫�[��mL4__l%koPi�?Ԋ�Ǻ���W���D�QdF�R��RG�eJK����00c�1�%9�d_��;N˸�edO.��ԼBZ)+:��%�q���t�QM�����0�np��!�ݝ���逑"%�ġ�$�CB�t��HKKw���|��p�;g�v���|��u��Qڷ.�����_���g 2�G��Tt���Cd�X��+��a2f��>)]�b�w�(�"$�r�����
�	����<}�j��8#��7��A�ah1�y��X�N��͛zomI�J~N�㐴���	��t�sNyݲ�`G�a�*����^���`t�0��������;�Ǧ��cu�љ�q����$:��w����!����]@�)�.����4�]x�����ӗ��(���|
4�����,�Qg���b��Ok������p�b�s	d��E�Pn2^�]*Y%��Ly(�z>=!��"��dO։��?00��`�U)�����;��z؎A>��&��I�%�R$��S&�ﺁ��})��U���kaW'Ĵ�$�f)�"�����	��#`	�a�\Cї�o����kA@2f�����et�KWEv�u���_L�B��.tm����~/eR��a�+���
�Ķ�/f&�a�`2;K
��0���%��7`�Fm���jk�O$.�{.?<y����b� ��	��i��o":���{9erQ8��$��Z>]�M ��/��	�_�I0V-��S�_d�A��C';�ʻ4:�o��u�V����z�e�=ۻ�$W��u�*�9[a��nrS��A\RpPs��M[eg�50��� �<��K��20)�n��*�#�V�B4@�'x|ɼu���ui��6l��5��+T���rPt:r��e@�@t&cB@��ҦL_����ї<l-�W��Y�l{��d�6V�a�e��*rî��~1|����	����D��z1f,��#�O�)��9g���+��5fJr�,kG�N��0���/i��W[A�_�i��Ѭ��梮��(��rfn��W���B��d��7("Q�������4����������O�~��)v����w.+AaϿS�2t����A�;���,��3P�uQJY\�����9������Z	�f�|-[���U<4ϜE����(��^��朤���,^W�z�f�\7���QN4�֯I&Z���z�T����z)�C�1v}Eҽa/Sh�kǤ�$�Wi��-	�Z���vk���T���	i<�z�<�{/-mZ8[��C�����}�H�j1Ə��q/��b��#嚫����L
�hJ�h������|V{��xs�#w2��s&�z��l6Q����_��3����\k(ٸ;�˓#�j%��{����^�(Y���[�e�<dJ�Y3��f� ��v2�K�2u,P`>� ��}$�"���?|��$LZъ3Af�!S�C�p�׽�Aډ�D`��עڵ�&ÿ[t��ͺ{o�����1,����{{+�VEݞ?;��ο��^P���k�
���d��?ߔ6����hc2�����'�mWazң���L�p�ճ�3�Qg����n��0�a��-����(�ö T[{w���hh�[Q��B执��N˳kY�q�H�����5�N�ĺ��Iϊu��:εd��\<���-�SBβx��z�xcr:����GD����yMڜՂ��J!AG�y
(q��#��)�7��[����$�Q���J��vv����]|�Gb�2��_ȔS��Mա�U=\TIL�<v{���e%�|���,�Ԫ� ��1�ė߈�0s�W�ś�x��������1�Po�*̵��mD�����<>��Az�E�/�Iq�6P�`��s�gۜ-��\ʨ�U�T�i)}�a��p�����ðY.������DU��A,]���t3�=����-=�Y鴃�o�ɵZ���Ib<}o��7<n#rИ�ٽ��vdD\��ձp 1Hُ,���zWx��C�I}�{h���@�M=Ǐ�G$@S:����z�v���ctW��EEp���|�*��(E��Y�m��̻����������1E���~`�L�ۡ�Q��P�lw��R���~Ppzv�Q�/]IW�3�d�a8)le����'z]:DR���:��>�,�f8l�E���.^�<��sya�bl^�[3��vG�|��-�[W�[�Չ �(�F�
Or,��)�@�*FHɔ�Q�L�_��#�_\؟0�o����2��Bw�������C���@�&v?b�6$��m���g�Ў�0Q�׵�����l��C�~�+�"�� ��uWww�T�y*�E���M��c�\��4����� eu�ّF��U/�˶Ҕ��#3��X�=zu�ᶮ/��N~BL/dU~5#�����5]>�T�lYtj�}
�*�!(�Zo���/4�-o��ҍ��Y��@�	���V����T�Љl<,�k�<���ΨbL��z!AR�z���GMe��q�Y7Ө��� ]�]��&%�p6ڜ$�����}|�I4��d�a�����i���aw7�q�P+��86��@�*rĦ�� ��֕�>���;�(�g����~ �%r�0����_|Q��|����E�d�\��cC��Z�X�F�;���y( Z��"��9���l.#'78>N.,<1{�)�&X�{Sf^�u��ٲ�� ���t��� �P.1}k�O�C���q��ww�l��蕛f�����f����G�&t��G	3[՞�S$��ēXk�,&u�%�@̓�%	���C�$�����gL�6�'C��'[�_��1t��k����T_�e ����a����:����������A�J����Q)������.��N�6���C�^�<J�ɐ����:�V�;�;��w_��_@@zZ:I�%��<q��4>�	T-����<m&�Z,�
Q\]�@��p'�J<�*+j���V���yS�B:��ڑ81D������?�d���,�^@�%M�q�p���-o����C���{t����86��͝07��� R��)�Wf��
�bҚ����LM��{�k�S#d��O��b�$l�77�[ �w�Í��b�E?N�}�V|�g��N�OMWm�.���3���Pcr�;S�b�YO�-�,fO�r���]3��N�"��/�U�E��e̡�͋;ߞ0ߔ������'���Ż/T+i�r��>�uӭB���O1��U���<#��[�W?��"��T[�+�dr]K���U����ء����[�wݳ��ӣ��}�V_M�%��>l*�8�x�RB�',GQ���?Q=�3��M���8fF� �~��`/h��}½����Vx�Q�Ʉy�D��ս�1[��'`c�J�0yҏ�e�3:�<�?��ڱ�.~����kА�dC���q� 唾�2~�Ẹ���"��v��G�v�Z]9Y�8Lb:�)�|K\����� 0�Hg-�	X��Ùt��m~���P_,��}��x�5�o������}�L��sK�>��NKT�wh=�K>6%ԺY�I�^�)�_�A�a���U�i��y�{<��K�
�(��U���60�Zm�957MJ�_577?xI�Y�t�ߣ>�`R�d%�Lx������]טt����7�Ψk��q&&՞�`	�8r��65]>\�N6b"�@Hs_ϥ�=���S���dX�4���x��O,���R�&�d+m���C�FC�ㆤp�,}�?[5��r��"���yb��7;Jd�Z>}ֺV���%��c��j��vv<%J�G�Z����Uo)f������7��Q���)q2����2!DW�q1���3w-"�Lr�ƾih��F*��`�轩�����Z�ND
���އE����'�K�*	�ʽ�`4n#����Ͽ� y�AO�hF0�J����_���,X��8L�:[��o��[|ȂW%�p�B$������X�4&�`�n�U	0�?���-)�����q�4��2��:�����q�\���䈐)ˍa��f1�6Ã4f2+�5{���ڨ Ln��+�:�e[���F�Re,ct5�U6ާpΛr�=#�_����s��������s����m�G?��yq�^���:-w�v�ey��҃4�O	�󹆝n�%R	Vz7�����?3���W]]'K�s�z\:*�1R��Ffj���7*[�r��=,7.��
J��c�z��������P&�_i�ty�Ċ9z&k������?lg���>������0B��:��u_�v�����T{[S�:�Oˢ"� ��fԳ*e�F��9�����T��j�ޗ�bϟq��0 �)X666�N���v�`�=�.4�u�S���R~jõ�1A6�"5D�bd�5�:�-M��[��1�<u�3�1n;!���Cgo2��5D�&�uߜ�+�%����?�jXN�	6G���]n�����f#n �\�p�+�CI����G P(��Z(D���2?N���if��~�ŝ�f���M�s�q�7���ή��ވ���hܙ���?�蚬Vo;b�#/�������,H_䲄���{�$����g���"�8!^�c��>��8��- �J����= �v��4�����[z<���v1'V���h�<�,g�'G���7�5�0w(ijzz�5� yb�����JN3�G�qܯ~�3�m[U(y�;*�2�V~�	�q�O�蚟Z
ў�v���xW��^�D���#h,޳x�(]M��f_N�	ѝV�s���M5�Ij����&Нq��vCSt�s]��{��*SZ��f��ZN-(L��Ҵ�2�Z�3�d�s�t�܊	�;<��&׻��uΌ�V��6i�=�6��P�U��*N;�2����a�m��⤲ֆ�Qc�|w�xDF~��x����y�s��)��m�MAȷĢ�٧�[�ﵮ6������9�<�&�c&\�:gy��M�;ch���;u9Oc�ޯĜ�\,ޯ�o�����n����m�����T.�6Ln8��{�If����ͶyA�7V�G���̢AB��yί��w&�|���o�ج��h������׳c�ZU�v1{l��*�f�*�h�ɯ��"��Tag˄N��,�I⾶M�¯d�i`I��h�G{�֮��Ml�o7� ��_�P\��CsAQ���:���Jr���)̙�ݸ)o(��8w�f�V~��)�o�~OaΫ𭸁_�}�.���Ӫ ^�+fd��~4�<�i���I��D��Ӳ����q }|�������ZW	�m�IT?�W�oom	��z4���+��uݴb½�u�8�)�� �_T�"ۅG�S5��h�t C�z��-�����$E��߭�a8���U\#G�dj�vYm��/Q�/C|�jgZ�u-�J~qe�#�%���9�Q3\��M�}�=��jҟ7/�R��G9YB����d�������=����/S+S���3��#;#Nq����/�>���}�?�� e݈���v#�H%�����"z%;֪���IT�IT�Z��o��F&l|�f�(%Uf�YE*Q+��P����6ep!	�q�n�TƋ�Z�)[7DR�I���8m�Q.�H���'�E��_�W��]�����5��)�p�ll��[E]�	��zk���V(��	��PY��Lק�n
0�tw:����)��[hq�z��*���ZԢj�N���Ԃ~mZ �H��)�j���-�v�.�S�Ɔ=:�Mu,����	�ˎ]�
DFȎRuT�}�F�9A�B=����l�Fdd�U7E��bl`I�����y=�d#�1G��.�s��ג�1�g8�=������_�D���?��/�6V�I��Û�Ɋ�q�U�DX_K�0}�&����V�x�~ۀR���_-�g�����j��>f�J�a���x���S4�p|I�ƚZ]{�C������#�9
B~-K���S7�q�ugg������4�- �]����#��ӎ�a@���O�����XR�yOC���{v�φ���6d:Nb1	���!J,���e���_�Wi��WW$�>��U��3�Pb�
�ǗoS�ܫ�6�Ve�%������ۓ�/GҬ/�;�Rg��9�@(g�)�{�0f0�&�R����;��J��9���V�����@X�5C��4(Sչ҇i�[X����+&�AϦH% E��C��q�>���K�{eM)D3�����o0��	�y���Y����V)2\�Z1�Y2ܔ(�������7�����4Gk����Fk�x�Q��"we����i��d�i �ȅ:t �.�7Y�:z\�rfG�>p8/���=�:�y�|��y����e��m���е��L��7�G/V�'凿}#f���R*}-!/�n���d�2cH����98"�k�@�x�/�"�羬��=��b�BĲ��
"-���`[/�"�xχ;���B������83��s�a<�T&�LG���x�F���y"	��Jg3
'�U�_�@���j���|:��َX{�����>�ߡ��ݦT���^SKj�=����ithXs��+�ЫH�$
�x��gdK�sq�h����e���R�!3sއ�l�����2^E��ή�:bT���ح�K�[�����؎�iQ�)V���ó�2��}�%-�T38Ǘ%� �Jp��_�i"ET�h��ϛj��#�7jW�I�)�����t�͗��TE5yV��_c`�3�W[��^d?vև����o��
����5%FF׫ܙ-�O��>0�ZU(��wo�EO����j�?�Av�m���"�上����l�7:y'b$pt�T�*V)���Iq�9�ahw���-?����?���j�xy�w��j�\�����خg[6��[��:�>yl��#�zf�T�ћ˧���k���y7��$~�P���["��U�-�}��ݭ�0d��1�b�aX���- ���^�yܥ�MB���I��o.D�$������n��o;t�R�v<�F�s��I���f{D�Xp������#�����$��A�)Ș%]O%�1J�W�^������
�pw?�3�b��
�?�{�e}��Rh��m�Dx�u
��L��;��|Z�4�u�Z�u��� �v�{B�R�/�\��/8L�%^�ߛ�;9��?���{Iqkƃ���#�MDV	j�}}G������������u�m�t�j�V���!i��[Aн��N��ח� ;� +���O�"�0k.?��%�M�m�q�w�q�_�еypX�w��.�����F��Ż��9�gs{�2l�7e��21w:=�b�	Ŝ�y/��,�au��y5#O�۲�}-ę����x�
J�ޱ�s5����ӂq����:��L���Z|���E��:�3���ꀎ8��>�� ij��.M7It/*�s|ѽ󉏔x9b�R�?�Y2ōd#())q�A+�pO�:)30%����SI#��]�vp3Yt�s�;0C�r��E�\���⌍�$r�س�������N�/��W��T�o�i�*����@c��a#U��
L�:�!*'���g�`11ߊ[�P���x:���8��ugM�'IEX3+��B�c?s42�>̮sk1�TI�e���z}\���}&�����!���w�sL���%e��_ӌ�}gfS�t�4��K��W��T���zKw*t$����ͩ?N1����g&Rqx���؉�����RU*�M�2�F2g ���e}D�;��������[����ad5�u}aa��c;�]ᾙ'�>��"[��FO�i�T����UKw��uK��)W8�E��<Da�D��i4����R�	�|�&�Aޏ�Z���^�n��S��}�X~)��]����U;s���ք������2��*��`���՝���5;RE�x^6YVx����5.DK�a�lf6޷�r�OR����y���XW��ʯ�����q�0��c Ćp�u��|�KY�d�#YU��z�#5�c.W�}ܘH9Ş(Ѿ_�t�j
��2��K��	�fuϧ�q��(&�1@������[|�fb:�G>�y�R�<?��1��kxe�r� Faa�
?��+����S0���J�|�\VBe%2& Tf�"�_���L@�ۨ�u�R���
~���=�7Nޞ��~���Mm�iհ[*���Â�#(��?@�9(��E���[�bYmfz�mn��E��u�� ��BvS<�H����O���.��_�?5A��!8�,!V�<ߙSO����U����L&�HQ��)���i�Pٲ"P%�n����w��X�ݪfNA5qr����(I8,}�܊��
n
��2�L���\l�̄�GyzE��:�f��8��>A�dX���͞
<rk�x8��"��&��r
R�Ц�~&�K�5S�״/�V����|=Kq2(C7*DLW���l�s���`#Q[��}��:�Z�jU������t����.#�=�>o����38��q���֨8�qx�N.�a����y�D���=��ϛ��F@�
����$�D9�Yf��?Ԇp��D�QV��P.�}u)�B���Ð��{�ۇ]��Ld�SϢ���[�|a�Gt+�DǗ�u/z�J7N��n
G	��[٨�8y��XdP�f�5#��AQ�?N;_D�]n<YD/_���&'�ն�� ��~[�����b�U��� �̎�;|fԠO+_MҪ]����I���Z����Y�~�����a]�KBV�`��f����#e��G�:jU��"�g�,��'�q��8��iR[>\�Q�.���ü�a��xS�!�Hr0j�������)�d~sl�;���
r�Æ nA�����И��\�B�ZL^.̯m���mQ�μU(�J�{-荈�l���m�Y�xF�l����N�l*1^� �X:qU�G����>� ��Q�Ȓ���r��vMsO��F��i��nXiJ#?�8+&�X&^��[��Ыnj�U�^z4�Dp;a�t3)�6�����<.���a������6d}@ �Z���E��H�g�6��2��n�oZ����{��	��3�ЯJ�	�sVa❿���b!RgC�����f6�f��AJy��`|��J�0���q�x�0�K��[9a7��5���_j�%v>%{`�}נKS�j;X��������Q;v&�v�{%��޵�e��@��=P�-�|�� ;��n�hc/V�r�;��,�Lm��ʰ��tC��m1��1�[l$D7!zӤ�qޫ���ī�͜�a� �opw��� ش��/�Y�}�]c��F�$���B.S�c�|n��k
W��Y�_���~v6:dD���|3�,OG5�:�w����KZ�����Ԫ��-�V�f `���H�rC���a���p��<�Ҷ�x�sqw��]o�^��S�eH��?⋕�ԨC�m�RQBF����\�\���L���fiW�'���)b���N�e?{+^�d��?V��R�-?�X�D
u_K'��3�'�� 3�]���$��V-	l����c�r�����2�cu�
�61�g��Otf:e޲�$����|Ã߁[������q|��9@-��7��W1��mR�GR'�A�:[%[���|�W
֡xhkM1�����9��7���j��CN�I;F�Ά�~�F�z���3��	�L�̏ȯ��YL�﷋;�[��s�� �'?�*��fiJr��i�7L9������M���Y���}�a�״cCgʔS�!l<Y����&��j�Z#^���d�R���|#[��Lb=�͜]$'f��m���w�_
��>��W+�Ps7T��x5?M<X8����������t�2f�]��0-�H������d6���)Q�&<4	f;t'5�$m=��An�
T�0l�F�����S�w���s��M��H|�f�[�t�
�l�S "7�8$� �IQ>�-�w7����	��ͥ��ِhP�\�P��̬�F��ۚ�x�o���3+��,�T-���N�~�י*g�9������K��*cT��蝠u1<n��b���x���y�����?8�d&�����y�o�+*�k���
�l����䳱����ڱg&�=�:6��ġ&7ςZ<���.^>1�1A���v�P��_*g-)�z�2e�̤2�4wr�A$P�;,h�W7���/0ʹ]�H�S��H�N��d���I�1�m_s'��?��k�'�U�,�`��1�δ
�&��+A#0�T�y�k�|#{H�>�۫(g���}k�Y	a�4�dh$`ѝ�(�Wx>r
�2�{]����$�/��O��سr��R���I�-Gq!�v��n���*�n��f���2c��4�&	;��B�1�s�;��H�]���oa�Vc�Ҡ�g@ҡS:�u=�`_��@S�<<^q�� �����<
��&���x(�����z��z�K[wG��4�	�~�����!:���x<e�l՝�2�D�nm��N'�T8�]�gPZ%�=鹢��u�[���aqj��J6���ѪvE94=�NHK#��7�������m}`�����k��)�������cU�quݜw��o�ǘ��V��K�r8e��.|1�14��4�����-8�Z���`]��<'���u�<���8�d���3��H�/SqÍ��)�7��Rtm9�-�WR�VD�Cz�߸��c�Z%ٓ�R1($,��-�`��lp���O��FP�!��������%r.�#���T(*�#���ILİ�^.�hD�W!���aXd^M����8)^gE��[�^\��������Eof��?֪`���2�M
/�T"rnjxxxn/d��7D�"�_�d*&�bH6�c�|�D���"'Ѫ�3�r����f�̂���x�?�~j��
�8Q��I������þ��֞[�x�W0V�O�l�tF��D�ͯ�.���K��#��1�']^�D�`h��J��[�-*&c+�ߏ����@�۪]U��&���ƪH�x����3L�� �0-5��MfL2�U^;6�S�*j
�Jg 9~��iW0�(&�� ���=d�/D�_�T���r�p���-p������cj��Jm/?�Z���'_<��6PW�(���R��=ya2!RUÚ��^u@���>�(�P���)\���t������OM��5��繓�$S��.k��d �G�4�Z�4�:��m��
v�b�z�JQ����r�9ik�:���?"d"���4c�E�f]�Қ���}����9�#����Բ����S!>�`e|w˿��RZg�L�(S]ï�4~��P�	�ɩY��]�N��Xn�ի+�(T_��H}Vc�_��XW$��)��od6�ۯ��AN��I��r�0V�><�R#�U�f3
���}�[��?0]d�L�f�z��e�:���捊�h�����{whU���?�Dl?-���Y^R��͋�W���݄�j
��}� 3m���(�w�ψ��6y�G�p1��(���J�H�~ K鮵���ZcA�����c �&�R!�y��HF�4���Rv?�6���F�uSְ�m��/���LA�}��U.L��S�I��L���Ne�Q54��Iނ�	�ٜ ���e+~s\�O���H�X�̪�\��/+P�m��`���E�-o��!����Ѷ8*���R�j��D�Wp@q$���,�@�<|�5�VY����g�?�:�1*�ʼ�rv��~4ϷƧ����tt,�n��K�aad�K�<�y�-?� r�r;Χ1S�w�V���]�zN��l�G̢#D�eɮ�?�W�"�>�x��OGtz��;�ώ���Q3�u^r�C�_R��$#'d����)h߳����-�Bձ=��/Hj}�l�ަ�hQj%.mR=>��J���%�����)4LV�*���9/��FUaXb�e��{B�s��7~�ī��]T��8��Pȳ+��!���]KxG� �3`�h������_h@@��p�G3��ۇ�D�I(���,S.:���&4!�}]L_�g��xް�9�Sp�.G��@E��u���)��?��w��7b�cI�5Թ1�
��}-��;L_�) i��|�/�C�b��d��=�t�9�����/�@�%�G��m�E$`�C��Xm�� tX��9���)���`��2c��h,<nƅ��(E�X���UC�����Qw�l�c�ޢ�>+ ��鑫�������4����O�I�Col7�@4)J��̹BG������FR�w�k3J�}%?�Q�����]��Ok���\b��OQ��1�-�S�$�Љ�^��*E���GY16y�xҜ>�Ҝ��Ik�ϖ�!Ґ`�`�/�zx��x3�zk�gy�l����)�P#�+�/. �xq`/��J�7|����#�n���]v�;3:��׳ɞ���)ad�� ���Y�>A��<X�8���q�튦8f1���	�l�&�f-��\ˎK�@��#�����}/H2Z��n�i��H���$5�'��-U�DqL�G�2?�S�2�?'ܗg�����m�s�/�b�����2�����fxU/띦����8��+ģ�8Q0���H��<.�g]\�(� ~��U�>`��T�.n��{��V%r�_׳�2�?��d'Ҙ�za�x��#���,�x*�ϥȾ��m�T�`�����yM�$� ��d���[��I�YX�4i ���9�J�b5E��� \�M�X��o�/����rw ����,�ӈq�Lޜ��(������I�?���rW���)�+�EEJ��1?�`Ȭ����j{t)��^<�?�)�l����y��s�A4�n[z��b�o�y��@5���+X���e���g��W�Q���OC������e��M�$#����f9Y��|���ꏬm�)5��옂�v�"�/9?T�7��B�t��	z�E(���~��
��?�����#*<����?B#y��7��n����-���ղ���W�nr*�7w65�.��21U�߀��h�������ǔ;��t�q֟
�z�#	F5S���i�y��*�z�a��=��ˉ���CʟT<�R��+{�e�q|�s�[ȻB�'Y������Z�����K�JBHMg�2��d:�&���I?=���=�������0��)��Ħ,K������0Ṣ��B���U���$�n���3�!�{���L���r�˟�l�����nA/�����@�7
�gbϢd��s��fw=Ȣ%�_��6�zn���0�#�������L���������𻅺��V�O��.�ك�U��e}�)�QiSrKۥ��9�?z�z�Z���*�p��5�u�t�3B+ۧ����H��I�v~uiV�^wC��~ꂌc��r}�6ɗɣ�n9V@�9�@Xr�6M�r>Ć4��m��珣�s0!=�� ɕB�_KB%M�DƬ�����7��Q���{Qo��F���Ly��Y�:�ɝc�����%���8�����.;��)���
��
*&n�hd*vxW���m�'�e�2}zd��T��lR+(�~������8��b<�&���������=ǡٺ�����~�&�� �c,w��Лz�#�1Qw,@�용a9Rk��C�5p���W���-8��\{��z�*��L΂/��c��ޛ�����|����W"å,BT =d"����ζ��D�x��j\A6��	�,8�_ݿ��y��C���Z��(y�y� �L=�$�&l�t��O�
�?b��)%*|�S�gװV챖�a&�!�{���?���t��V��(�s3��RR���Լ�ԕ�X�K�!^�ll�o�M����(���}�*O���H�抬HTFZ�hNڹ�up�X�N���}�r�.�WH�6V6⦉�)f>p�62했�k�12�2,�=����{�+�E�V;�֏�R��8ͥ`7ii��&��W0t��eP5���[���&�94��H(9 ��zX2��3���tumV�0]�q9Q�C ��觚���.�,��A���T��G^x�q�>{ø�J�ߚbz>�����|ށ�-i(���w)����;u?!�[���T��W��-�(<j*�i*F��F����E����&-�h��˫�|uCSh�W>TuJ��Pi���9�T�vu��o�X��\�v���
��K�����"�����CH
+ٽ,dL��3�+a���� �
��)�u�69A�ί髅g�F�N�
��bS}waceLb[�l�FVl3��*Zҙ�;��^/^/�|���/E=���E�fn�w��\߲�E#m_p��lJe��_���<����_`������ʹ��eB9�);+UE?��P��}��� �s�D��g��YP*	$na�d�:.�P���H�{Q4t�'
�Fv�0����e"t���h��矊5�+���'�BLn����;���`�T*��$i�:oL�������;�ԥ��9S�VY�����Nfr�FU����-@�x�q�Zy��{A{��l��u��('�r��Cn{{-��{�B �v$dD\�F��K�I;T�:3��oN�?�{���P1������0���C3���3����ϡU�%C�u�A�_�t(�Ԝ���&7h]��(��pM�/�;��o�^�B;�����,���Y�[�� x�W������""���\�cC��l���<)��4t��J�*�y����d���D�� a�
e�d�u(|5��
��u������raloq��7\ڽ!�� *DY��96X`b��\����@��Q	�A���]���N��?G�L>�x6�jKUCI<%��}�ia�������/XBņ����"�����+T��fV��ۤ531�ٯ_4^��7�]((fjZ�`�� ��o1��/��Ct+i���k�&"zA���b�L
B��Bi.��i���?��T��i�]UP#����1�Z@��_���i�����x|П��X`?[p�*��Ņ
�v(%�����i~�I��*�DGO����<��9�^��ݤ�a��I����A� �X�P
�w>��VN���p�>��:δ\����FP=i�!�c���BP@ �Z;����y�y^ۡ	j�ͨ<Z��x�Q�3��vZH�	�rF@���4l��`D6�#��9���<\<���
"�|���J�������-_,@��k���	.&B�hq��#��B:��� z�h�������G,�.%�bD��3w�x~I�8C1����%���W���I�\�����O{'K�[},~��;M(�J�9�&?��*� �P�V"}\m-ʏP����Q	M����-<:������qC�Ly�U{�	}��E�����,�^f)Ͽ��	���.�e<.����V)T����H�ۙ
�g�
U��o�ԟ�(�`�|��ߟ��5z�a8�������
RJ,���}��zΛ,�����W�!�,e��[l�|�M4�5j�'E���%yW!=�~�C��!�7��:;{�)g�&�I�;&�*���Q�=iX���O���˜��15Ǻo�8|6��d��}w����=$�z�����̮)H���A����¤��JUI#g�'�\P��6��)��N&�a����O�gZ����/4�[y��ÿD���d�>�ʖ�ozTP�@�Q�	[N8��6
�(�r�)�(�TA��Ȱ@�&+\ƻ��� gӕ�����e�b���rkj}Қ��(�e�/0��5h[')���ϸ��Q)޶���ax���$;��k9����*+��/�8N�����E�RQDG&�_9���[`齹/U�	V1L���(8��8����Y4s� τ��l-_�ݩ�`B*բ�L5G��Q��並���DzU�5�Ep��-IzvgP�j*ĩ�_�w��\�!�����Z��"a���U�~�+L<G��_E�#�@5�"�x"̟J��}G��N�O��2z$g�,�%���s/�]���H�(�a^�,)�%2,L!?�̭��� �� L��:i�;4��4�1��Pۮ��cQ�b1h�~�� ���C���2#Ю�{zJ�(
��y�4OV��Г9�Y����j�i�C�(�����������.Szq����&F�mW�<��ha���ΈSh����1�$�}�Y%�&]��WpR�|���0�Ͷ9[�3��*jͷ^T��q��Z��9��	��&�Y��������	�s���7=_�6e8K=��z"dV����[��ɳj!Tp6���ǏI,}}}�f�9��u��Ԥh�:1*,�Fq�!�g���>���=�X�,GN��5��!�|�7�Km�d�����^��y���#p�^|;�������,�@,_�	٫�L�mf
���O_�t�?���a�m礛"�T>�B��ps�K�#�k��yTo@Z��3����.O͢�<���W��%ۧ�ʹy?�!��Gk��M��"�T'k~)��
Κx�+��e�m�.���Fi(�����nݩf222KGG4���9y���SWR[݋�Cғ���9KT�����ӳ���%�eK�����]�*vݧ��3��ҕ���خ\�/:��U�4SF}��r�)�x�>�g��/��#��~��s�7L|'��do4Ȯ�w�d!�ǰ䤤0C���1xV˖F2f�d�<vh^��q�`2��#鬣���8Nw;�q����#D��Pj��JwJ+-�-=p�Db(�;D$"���� ��������gg�{���z����3�z��XI�>K�𷆾}�Ej>��F��=����9}���ʯ�Yh�P�S�{�?An<�,�'±~	���[F��'��W�t������>��w�d�p��{�Q��F���u,ޕོ����w`؍r)eT-A�ǟ����@��LQ������9[r�6�x=��H	�t1�Z���b�*Ѐة�F���wgU!��8�����C8��vے���e�߰ovn��l��)߀=1�|��Py8iHZ̵�*�쥎�ħ
1�Tl���b�֯Uc\f�+=�B�v�LIq�����oH�o��_~h~ko-_�?L[z��Ad��+�<��{k��!�Գ�w��#�Y�/�<ma�ĥ$���5x߮�a٫��D'��-ߛ��C_�2Ϧ�h��R����;�pxmFds�yԺ�Բ�G�v�i8��͏(b��W�C���X���Z�ΡJ,�����7�H��"%�c*b*�.��4����/#k��Se]�&�-@H���F��{sċ1F����q8� �K�Za�&�-+@*Ь� ���Z��$O�X=7 SCZJ~�@���>o�x���T���+�pU��#<�p�5���':�Pέ��W�gg�DQ
�b�] iضkd�iMHR�;Mb��$�=H�pMj6Y+�����ҹeg�L�N��A�1+$֖�1�4$���	pn?��;Tǎ*���Ůب��r�"S\�dY^�?T�� ���3���4TONɱgu	>U�vد�u���}�|{�.Dc)e��`�G� �9�_�Zݳ8}��q�b�~q�n���o-+u�����Y�>��D��=�8y��MQ��D-�ֻVQ�Z����h�ޯ��3��t�ܛ�|�SZI�n��it�F%W����PҎ��b��l�=����cJ�s�{�e����*���!v-LJ��|���>��l���c.27ߕb+݈X�A+�d��J������c��&�g�|Ʊ�pr�����!sǉ�
�%q��~�48|�-�M0,�E��ŏ�

Ӑ�s)���)Z�t ��.����/�/q�ƀ{1�s���h1o�d��19�����i��&�.Fs�}ڤ$'d�Fi�Ŏ�6}5)�r<$��@�=FK�Ȁ�F�4��C(˃%n#o�f�Hb�gm!�M��05���#]< K����u���O�x��i�6���0��5=�TAZO8��3C߃��9��-jRhbv��LJ ��b�u�!�Zأ|��x*��D��Y
�"��TǷ_��2*�m�#���y�f�Ll`,_ZD�s�`�頺��"��W,��&�sSK��]=���Uz����_P��x�?$$&�X�a�o��҂�#���,w�������t��}S�ʻ۹c��ν�ݢg���d\��6�1e
�����c�#u��������[���z�\j�s��� ];��{6^���H[�S�J�ڌ���#��v���:�i���6g�1 �I)a�$�A�N���B!")��ǗD��4)'��@y T�G0=/���Y�T=�_�2`N���(탊����g[��U�m�V��N�#oF������eJd �
�Zu����c|���vC6�K0m��R=�V���r�����%]F^�]�Cl5�8+��iӧo������ŧ�pn}#\�������#�Ȏ{�Ј�4����Wc'%P�^2xd�Q���i�r�X��I^k���D���r�����T��G5p�(E�W���aWs:�B�OZ��	�o�S�I�1;;Q�ׂ���*((45�B	f4�$����=����J���#���:4sXg8�4O�_X��c�	p��Cq�l��4�㌢I1�<��`oRf�/���Nq��̇��~6���6�@Bd���l���;�ŒD�o u�E�1��`NVKEೋ�1F��ɠV�����0�*����qL�$��<�ӏ�r|,g�|%��}���L��K��x��j��{*l�BiD'������1���cu[!8 ��Z�����
u����ӧɸ�3��H�|m�7���CLg�p�e:�f�IB��ݑ=�V�`�M��CZQQ�������2)u��7�Io�c�0�Ri���O,`���|�'|n�r/���Q�u��� �Uʛ����=��اt�ɒv���W�9�3�����m=������W����76��j�9��9O-�?Ns��c[��D���^b�P�3�뇍���$bcAt���Kg��/?���/Z�<G�ie]��ꏧ!���L?���h���!�r�36al�^�:F��em�!l��V��V�z~�ֈ��>��l��=����[�/Q���x!M��-���ya��Y����uЯLN�e��f�3�]���K���1L䎅?��$�yE^*D�a��"C����q���P"��JO�V�ܑ٣j��	��K�}��������*��?�6�}��r-�J&
��V��f��,��!�u:�LYV�C���s�*l3���K@3��݉W=;��^��K����7�X��K7���݅&d��+k����(S��z�>����i$SG�|��޽�k^�n�Vk7A�(>�<��=��{Zؠ�QXR6-�S�̴@�9����X��~E����=�f|L��(�@�wp�ʎ�/k�����,�ƳfgTf}��n�q8��߳i�,����~����7e���I:O����8�}��!�Jz��#��Z�@��̤�W&���g��@�o�Q�-'��~�pG-8�������]�[4Rv�Η�:�jEp�$1��ض�;#��o��@�&,P�h��t��z�6�k;�>ä��	� D��B��N�7��R=�`10� �tjK~�zJwAo�ӄC�����6U3���,��������<�wA��V��3K��c��tpK��l�=��
����� =o�lG�ʂl��D��%
�O7�0@�J��f�L��l�����Q���ѷ�G��|�II5�?A�6�f�0����wN��JoP@��hE~��B��2����8��Y����?�ts����Ȁ$�Yc�x��>{Ȇ�rG���<������.T�{��9%K<JG�B#a|�1bQ0��>��纄�!���둎�[���+�6�m��V���ճ����O�T�$&�]o-=�7@���G��KH���/���w:k졜� Rf�i��i�줡��j�7��]k�)LA��"�P[d`K�U�2>�S�Uu5����;��3Pj�)H��de��芽� �{���|.�$�7Q��Wn&��٩?�nv/��a��AOTC�t�;�Pm ����o3eK�B7X������ǭ��$��0u�qE��⏼�k�t��,8K�,Vh��0G�JTTRrq7��V��3}���P�P�뉰���j�N�lOF����'RW���B��������Xp
�--����F{�=L�9�i� 2D�We���
��ϫ�Oz�b��cC&�����?���/��t�2�=������i�QyF4��I6~S�h	G]ʉJ�,J�G�O�v�~g�F�7�|������ڀ�-Lr�-�^;�D_~5�N�%(<"�M��ˠ����&��!�����pM@׻9Rz��~�s4�[m*Y��?���L���s�ߒ�̪X
&ѯC����6�@Ȓ$�j7,KO�}�7��b����yE�1R�����ٍ ��M5�*�D�t�!yYd����&���&�*�h�rr��������Tb�O�4�����;%V�ku�k�.Z�a(��Z?Bd3�?��>��%<@OX='��P�̠��q�a��1B�'lb�{UȠ,�£9��)#�4�ɩ�uB��a���) 2n�Q�V$�9��߅ ��m���d)�5�Ϟ�M'�J`MQ�Jb~kgөl�@԰�o�,�ˤ;4�(�S��=v�(��xf��M��pbho���-}�����K߈��C
O���[Y����Л���ʎ�q0 _����	Cj�)R�4�(��6wt�����4fw���7����+��|&��-�2�N61����o�/��/߸#>v��d���xJ�Vw�#�f\	��e�ܨH��B���Ù*�^\�@X�� Ɠ7��e��b��T�HWD����>��{k��^�*\������D(�����1A��eG[NLTʥj\H�e�GZ�v.1q�f�	4���qg���8i��k-K��LX(r`0��x���w8cyv���)<h<�����h,Ƈ�EsApsQ���wt�Vu���{�y��ğ�l�r�/'|0��hQ���̾2o�*��b?��3�xpט� 1��4CI�$~�@�ѷf�Pz�>��|�[��yXs ��,q�}�7N;�	/�e!��$r�ޒ�ƕ$JQ��fgH��V���	(d��\��]i;4������+w�k*r\�9�a�xg��q1�hd���nN�\����KU�%VWd<$ɞ�
������՝��qQn�}E�S^�����$v��Q�鬗����$����ٍ���z�6�d'RͶr����rq��������Q�k�hu:mN��hj�Cj�a|��v-=�7ݓgE�ZF:�ׂ�U߿/�Is��b5	��(��l �C�@H7���E���f�7�<d�n�P7fsIB뻧��c��>�+[��м~Ac"a=NC���\t���@*dV)���8����	�h����v$9���z�7�(�@Uo0�y�Ad潼uN��{��-h�A8�3��tc��C(����R��|��%�R�3\�/:-��׷�0V�̜	������@�Ot<�]Rb*UN��s�xx�;5Yi� Q׀��˙cx��,q�fH�f*[x�_��D	�O˱P����y:m@�A�6T�&���]"s ��d&23ۛ'��,��(q��͒J�x-ANNNbƈ߽ kx��k�$Q҈�yV~��؜��AO���X���my�[�w��7~yy�ܢ5Sh.�*Y���Ջq���kZ�i��I�>�b2�y ���i������4���]��^������oiMI~-�Tr�+�8a���ݛZ�7����4�?Y)0D>�e4�V�1�����d�c��g���e[O/��_!���.^nj�E��>�\L	6�oe�-�hM�^��6S��s���ͫzic,���Xz���, =���+p�X$��g���[B�9��j[�Hy�=O��=�>�h��̷�NrJ��e>��Ryf�48�ș����:X6�-�%⫛��\Z8� ��aŅh��*�ٜ��x}��`J��&RR%S��Iu�����~F��wW���MK0�(��X�=Z���pSRVl��ܜ,S���+�_�1�������)���Tå*9���mSsЧ'�Y9@��EY�qͱ
{�����Ԛi5luN���r�r=S����l
����L?Y�*^���)-��;�J�q�@�E�]M?)�����Y��9���f�K�i�ʨX�e"��C�&6.�>@�S�veW��y�1%�A��ȫ���Y�d�������?�y������I��=����x��H�C�'??S&�X�U2wI�DAQ���!*[L@���s�T��Ym���e���9ir6��|d�9!1RGO~���iN�S�x�G^�+��"�TX��Mʉ��@�D��:����vh��N-=�:�ȣ�a
&ePV�O�c��p
Di�\W',P(ٱ�Y7�kn�_�������P%�g�L��_�^�J��N�X(�X)H�Bɿ���Hl�D�Ϻ��q<{�ث�ӭ`5�}����@�f�AG�������������D�9>opuumjj*�4@����l���m=��zR[��:#�
^W4j�y�A��!:N�)��]n'rhn5�.n:gl^o2��C�b1��v�ߓ+B��x�۩���];��N-P�S#Ay.ǎW�!s�l8�D������F��B��&���j��2?t����aiD���ҫL'�x���S��kn����J��1L�^gʏ��%-P��H�C����ԇ����ok����3��2�:�;�S�膘,����&)��y��O/�}�u'����.U�^��F����9��X���%돐�/�J�ļ�D��p���ɨZ9a�;v��)��&M,���g��y�f�CH�uX(ft�q3��a���i��cW!��6^�l�:�l�B��!�����4�ż|y�R�L�P�K���]- ��	K�����ɏb���	Z��绤��P��.x}�J�DՖgrh��xCͶ���b���d
�TrK@�6������&�=�"�
����q�x�!oʿ���zNcT���9��k�����::3	�f��PQ�e�.<�n��f3h?���q�Y���.�R�5�l<1�L�#�4#�})@��,c%�gB�,/�?�J�^��F�Ě7Fc%*��i�S�G�9(��_k]���� ^�kaN�3h���r���k�f�9����]��y!{������1.�Uz|���df�Yk�-$��UF"�,���Z:��[��Ҿ��+
����\y�k 9�ct�d?J���A�����J2��:o���~a%�����3'|�ԃ�zD����L�|\ϡ�E=�w�szӧ��t
��[�����[�C���6,&ĕx[�Q";�5t���/��K��C�-~`Cr22�(o��}��3y��Y��T`�~�7����0���Ok�����32��O�����,a�2m=���dLkŶ댐�+���(4������6Rw�C?�c`�5%�E5QN�ߧړ�����җDj���/:.N��X�9��LV�Nz� +¿����@%�[�ѻ�3��S�VkWiu�h�8��d�ʋL�n��q���Ө-���L��<�Y�^�&�Y 5M���"D��:j���<�̟�3�.�s��]�^����(��l�J^ �?N�k�.���C�@�B�����)��ξN~c���ODW[7���+ӻ
�ވD�<��X��wNM�?K�\q��F_Ff���9��D�s%�p����pl����E��C������j?<&@(4���2ţ2��HѦ+��ȟ�	J�
������%3��g���ߐ-J&3��0����C�M�SXfᷛ�X�9h��d�!�I��jG^�D	�������9j���q������������v�TJ�P�+Sӥ�8F���|�vUqMkυq�-�H�;;��M�TMr,(,���u�q뿵�����o(\�[F+�EG��$MۑJI���ib�<����\:0�"�����!�/ �}�x��	P���7�F�2p���cu�-fj}�l��{/^�4��mĹ[�@Sn�\�W���?��c2&�h�43X��ǕT�����Zo�x{�Kڟ::$�2*jJ���9���gvOBO�C�s��ribI��\�gMĀ՞Q��}R�zD���cj4�j�2�'~:a9�G%���f��r�H5�g&@Ctt��Ě��돌��ӥTW�f��k�_:=����z�O��;�ZE�{B��G���"�YJ�
��W����G�擄��78۷,,��pJ3z7�4�I�՘i�>���B��:Ix��M6��0�Of��ϴ鍁;^J}���K�Y9)�?<6�.-C�R7�{���~��� |��Fy6n�m�l��XX�جW<�t�i7�>�mwe
!y����}r���Nhd�u{.H7��[���V���W1�n?ǃW�� ���]�f&xfm�O�gs:(}��ʏ�v�c��k�7��5oi_Eh��n}�[�t��k��Z�r�����S�X��c:�=|)y�5���J��8oĥ��F¥@���-��;ʵ��ZrgX/J�J.�[�����!�䃔���1
v���3\Wh�%7գ�Iv8�eߌ=������A�ɤP�W���h���)"�r�2�"��<��U�~l�E5|-z���������qB�K>ۗ9���<�Ac�?��G��422����~q&��A@Z0�L���!�]]����gx��E�?���W� S��n=F�5n�i��Db0`���(
ӱ=j��).ml����9㓁Ӂi�%O%�������<�{fճ��7W�N�'���D�Q��WׂK���e��Q�:���}cF�s{D��Y��']%#F�2;ϰB�޽����s9�0X̸[D4��LҠ)���=y�"#�GtbB3��bzJ��/�t�9 X	ǳ��uy��L���;ͻ���&��7&��F��=��eu���/�%����3%QH� X{�,v�mJ�_nF1����o�~~S[�<?�I�Q�
��Ix�"���DG��I��R������ID�Nя�����T��7i�*%�l��^��I�>`G:�85*�1A�y{/��!���Ynh���d|����[�����S�R.(MP��@ڮb��H{�BҍZ+ob\��g+ƀ�u1y� �N'2X�� ;n���S�.�"ϊ�+�q�F�y���Q��Q[�����&
���aA)�CH,��w&@�	?'1 Mx�MR�ڄ�ɠ?����*�;-���p@�6�m?M�J���:x����h� `�.�Go߾]��_}&���#g��ϲ��ROŠ��~;L�m q���DLZ���m��`�K;w�Ƀ���)���m6�hP�W��zo�n+�(�:(���%g���4L��{Wx������bV��)��K;;L��y�n��w�崍7_��Q�e���@���f2)@��naN�tB�'°��vT�� ���Xe>��[K��e���\�o6ڰ>%� U�[�`By�"�ϥM����N)��U�̩p��S}��H���ۙ��]!��[5h�TO Y�~��9#�[�1`��k����r��IZ�SS�1R�������b���a!�ڹm���ӭ�Z�FD�hJH�������*�l�J�!e��^�R�KpXmO�o�;t��O�-2� �L�a����t�}�l�������yķ���,0����Dώ����C��"vfr
�u�҃Q�t"D1BUPG���[���j���Z�;l�r]/�;J��޼���9��}��t�FQ�-��&6�6>�M4��jqռı���H���'1!B�tГ?@|
�#�!Q���R"��>(:�>G�kU���&���_���ϕ+z�l�m7�/.��>�J2NOO�͓�����d��j�V/y)W58�@��Ĕ�u��e�ӷ�/1X�������j-Kܭ�+L�fwO�*S�̢���A��CMMm~{��ZF�9��*������!+�t���q�IF������o�&m�=�C�*u�o�G�4���v�A$)�+J'bt����I^�aݕ_N��i�w"�=�����̪_�^�㿌������c���5�ik��|�_��2+���x���L��`�׹U�`�6����4P�w�U�r-Z�Q;gm�m[��
`�w{�ڻ�+�8�阷�����ųBcul�Q�����%d&y�;/Ӿ�	e��ܭ�U�@�2���Pɜ�hݥ9b���X�Ʒ����U/g�h��؋R���agN@>�1^+�@g�m~k��;/�=_��7�q�,	��^�����˽����s8��w�q;��&M������AA131;_qECr|�2?��e�Y�	����hY��̠P�Ya�яic.13��*��y�%WU���at��(����sޱCs](��|����(齒D:��	*�cR�i����]5��{��%/4�f:S+�G�j9`n8\U���1����7����/!�\���Ք�=h��g!<����KnuHPa�؋��J�KK�t�ƝѠ�n�v|k�OH=�i�����^�5��9a=Y����ꔑ�����s��� �l�5���w�<jU'���	��B��I��l��"�?��D��F�j�>=cs����Ot{��[0`��^���ǂ�7���pyO۫��0�~�U?ΈJʈ:��̕W����{��{���f�����b��W�?qj����ɗ��Q�Ww��1����7GIR��"��C԰3��ρ�G���/�wT���y��IB@�`"�����!>=t'�K1�z4`A�~#�my��� K+��/�s)rQ&x�Ĕ@�R���GY�]�.�a6���U�8�S�9����BޞVT�����Wh�UN�Z:0�+@��8P��|�c�r�-���.!wd3���xip��t���QY�5P/���r:�8�6TC�h����:ع���~r��w�8*���-X+E�1٣�aƍ��.{����ǵ��gAo=�|����y_i�K��hU�?���M,\���qN�QG����ݛz�T�g��Y���e��'x�-_߁o�Kg%uW�e9qۅ'/��*��֋�A���^=چ�aN��$��1��yV����`@�t��\=N+Dz� �Z�m��ne�ħlCw���S���W�c"�s1t�p�@wلh��c��Ҋ�	�
�Ӎ�6��/I`�J<d�I{��B��5�4�6H{��;�TL{e�͊��(Gd:��;yJJ��d�	GUR�څ��}�ynhK�̒��&C�9C�z�S��F�,<$�?1��6ә�{G��a��Aj��n�ŗ�ė\�Z^�jW\���**0S����Q���P(�{u{n�~��������7B�����@>j����ͣG�K1��/�v��u(2�(�
�o�x��A��YXڿ�,雘j��a�薖�U�EEO>6�*��w�JU��]ee0K�p6P =ߢ�ặ��l���%���X�G��$�z(UM{&����i	��9~|Z2�z��=1�-x��Ft�����v�"ε��</��^�is��P��R�� �^�������=���mS	��u��L��ѫ5�����+�LgƲq@����sf�����@�<}8`p0]�P��L+�/���~��{M19T����麌}B�E��Q-s�Ђkd�l����e�P���w�b���3�'D5�Ia*������H����|�y�G���瑶��#T�>K++��B�O��s�ـp�P�J�;�m`OK�P�F�^��cI�x��N7_�a�<K߳���5M��I�͎�d�N]|��E��@��	}Y�_�8�����>n���&�γ�ȿN.��$:)s��琂��.��c�I�!:����B�cg]�Zc"4���DR"14Ӑ�㓌�ׯ�G�r��L�Y�=���<5��Z�k]ܜ�kN�-Xj/2|uv��a��c�d6v6�7�����G�@rp���K��3v4\�}�.�VL����7�`�jW�XJ!H���N���/�"�c�ѿ	q�����6vvvn��]W�A���R��2E���q�=�ъ����fm�T%.��iKzf�J��t��BS`�g�=��s߀��������@Ư�,
(��*rjƍ����t[����x�x���}�b��#ѥU��5 �.۳����}��g���t	U�d(�!ؑ�����f������'���}��ԩ�x�AP_�_X�7/g��$��cd6�f���~�K��l5_akMb?A���1�C�Հ|��!���^;��ZA�@�ƌ�L���>yF�yk훐�)� ����M��'�AAAa�*3���N���6��t;ר�x��1�$�CԺ͟$�߶&q"f��� �z&�K+%-�0{c+�g'�יj7]�#<�p���i:=P��O�&D],�4Fn6��^�_s��[s�)��{.�|w�J�?�P	��u�t�n��v����r����]&j62�.�{��b%S\W��O�Y+�*(A>J�^�iC�g��Ӕ.nY�^����梜_��/��Tn*閨��ם�NB(�ݬ��H��.�ҥ��E�
\����{ɕAJ���������)� Z��uV~m��-I:`�N,hO+8/�ȏn����TX�E�f�ܤ�&?�{;v���vZ��r�$� �n�J���1�q���O���ʹxI�^�*�Y������B���~���m`@$��֠�u�X8�q��o��,Ϲ�W�_B;���!zH�k"V�c�Q���� ��=e�ݎ��'s�~��37�uAH.V�x��P�L #���g�&1v�������<$H���%E�D;��O���U�EA�ǁ��i"��_��]�F��_�.[��1�۟�|ga!����G|��Cc>�i"Q9X����^3n���Tf��=ť��[�o+l��{,j3�P�#Cfk1.������W��c��f���������1,k��i��_�Z�W��Y�����[�s�\�� >�*/2�e�Wǰޒq� h�5�,>̤��.��l��lA�N9}�-�6�j3>��ʬ�
�JL�>T��ag��;��6�&���fwwB��]�T��]5�od�v0���$&u	�z��o%�!�g�VW��NI:$g<���
ۑ�=JR��$�D<]�U����ܬݼ��4 ����3��ܪ�.%;�'�_Jk��:�8���M���ETz,1�r����;��e����}�����}�b���WeV"G���"����:���y��r�6�+�W�U�:���'�.ī�o�#�y9œcqo�%y���āo��|].@b�����9$��J	j�����E�ĉ�,��)S�j���M�W�*��;��Α����g	����B�9�6����7��z+�oK� � ��Bϰ[C�o43Q=����|F� 穪�p(i�^�s��C�"�`���7m� vH#��o���ث�^���Ӊ�}}���̝i��~9�s�u�X�g�����H���^�����9��͔��8di1��`u-Z?�\�w��E��ƇGǵ�`p�콾f5�>{Xt0;����+)�!�P+��r�?4F�^�����ôLԬ�o�q^c7��^\Q����L��U�_5G�0mR��MEnv�t��8 DEq���4~[�8�_&l<���{��s�g�ڄ�1��4%��)z���+�K�O'˙&�fu�uɏd���4E��woM�u�ķ�&i�Y�ߑ�OY�}��A�=�%i��|�5^�����[�C�������@��W�ރD�:����{2`)���&����H�(x�*�Ѭ6	X�`�Ƅ��@�c�"�d �kad%	0�.�lp��U���s���WS�r������ၩ="g����/�!AiXo�wo=��[���Au��x��A:��m�eF�/3Tj;��D�e����T�lE���p�������eG������������,��������d�ռ޽j��?� �ڣ������?qE���c�yȓ��2�A�e� �ꠣ��j�x�lz�_��Ұ�]K�]����� (mh���k&*7�c�	��T��Ǡ�18��@Q�Q̉�'��.�3e�����c4���,8����A��;M����V*�1�A��}�F�Պ����3)Yƴ���=Q�T'�rdRK�F5�X�m���M����xod�&�=����'&� �D6�2�@����Y�����w�9c��������ݦ�g�7GضN���]6K<	KC��8~���7C��n�P��z��b�^�x-��o�DP�p�p[��f	�G9���H#e���Ώ�;��2�aG��p�~�yb���vX�А�x�kQE��a%9.���ٌ�@�I]�y]Lb�f�]�!��LP�� ��D��*���ʮ��ZT���r�m���GX��9���o�-���5��4j�7�����JE�~Q!	�,{)������gy��o�˨Eh����ҩ��+�;V,P'��A�=�%�����5���̳�9��� =�9Ų��)OLf�(P�M�[���F�O��'ug�o���w���4���8_�K�wg.h���<��k���s����(��q���Ape���Q��S���*���M��5��O�l31i\�R�oOҤ	�})��h��K�^M�b��Q�!ꇗ����E�Rݶo�ޘ�i�TZ��B#�G�Βi��ɒ��ؙ�ޠ��]��0B:4�"ʊx�u��lS��9¶.9Q�4��؃���v!_%4�)z��5�����I	J�ڿsEyu�v�n���0��TO���.t�(�֛zN�T��������uA3+2Y�����o��S"��h��l��x ;E�s��R�@o'X�#�[�(l��H�z]9;��g ?��$��BT\5��w�ļ�m��%K�[K|�ؖз
���mX�8e��!iԉ�C�8�&�i<�>!Ln�J���xh@�evo���I�c��.5�q���O�t�`,�!o}/��p��.�=�¬h�xW�+�w�ty�.և�����,}l�|��ڰ9��@����}�l��'�Âϸ�vz�P��C���XHZf������2��Β�u+%8#B>*�z%E�5��m�s4b��a�M���=&h�6�z��W)���R|�B� �i�0#��l�9�B[F?����#�Н�]��A�_�.�0{������=���ژ�S����fC�<�^ �i����_��O2�N/w#��ko��G��;O�N��Ĺ9��ɾ7�9�1B��b����96{������HJ�3";�	�n} �:�3�3b��)V�0�������7n��QUy��ھ���%�/�� �����Oq�"���	��8܏[$U�	�|�~P���'� ��	�W��zO��|��>����{z�A�p4N±�9�HY�;h�X��e`��k�ּ���?�g|�L�@�Ҵ5��[b�e���դ�v��jtx����|�겊Yt7��^�9�%��ҩ�2�u	GP���68�R��C�0@�t�qpC�,��!D�|�F������z�W7������77�D�y��\<��+M��H�<<���w�mRE�y���TZv�@����1��=e:cA�(��p[��i�����z�p��ʏw��w�̙I�Z�մ_�G��F�
^\md\�����Z3�bP~�����AI�]P�YT�{��d?��^�|y3RwӖ}``@7���}K�����b��F~�e�������U��-${k�7�Tc1/��糙�J�%B��IB�P�,�w뙆>�vd�&
(F�������yϐ\5p	��cw��l�\�|,K�\h�}��k�l�Y�*'Q��,�E���:��4�I0��e�-vʏe�1�[���GcV�+�%|Q����Xm�3`YQ><*/!�Rs��|�AY`�`�: ���6�od�8�Z����3��:z[�5Г��~	�!�� p>�,��9| 6�8ÿ^�R�*��kQ�^F�E��GZ�餩㱉1�&��Y�FN��0��Mh D���0�𼹚�R���ri.�s�A������߻�Z��Hi0��[��X��u"����i�@k�u�\�]4V�e�\s �q~]�e�(wg@�׸{�R VW�o��
�X��}G۞�����E�v���]�=��K�-��eۨ��mĚ�f\՘�������i�l�d�]�,��p��X�>6Z�0�J��QH\��u�u�����A{dm?�P�45���#C��j��q)]�ֽ˄x��lu�}|uEb#>�z;O�J�T!�l8<��eN��"���c���p���2����	��A{���-��dM�;p@)�-�4O��EN��n0{	Z|L�q]1�ɧ���[�6��B	\��/�?���~����S�m�������@YY�������g��0V��-$��v��)w�K���{(�{ݓg���S���H���ݮ�t�\�]Ҍ��Vf�W�'D��%��0�-R���k�rX�f>�։�?��T��Eo�g&�>��3�a)��ooKݓ����'_��⢢�����2t����q'�Ŷ�s-��.0i����Z_��_ŝA����'y�*��ڊ�T5���4����)�D��}�	G$�F=M���{�4Y'�K���~O�K}����RpM."�u��^Y��'W�=��SvH���ꔎӔ������S�<�BH�잡.:s��	;�L�O[���|�������Gozk��.�#Y��Y��r����_/N�oex�#뾧���9}o*�1�Rb�M��V��=բ���պ�nS#Q{�Ǟ�+)w΄,:�����v#CBB@�t(g{E>��V�����R����@��sH�W=ɋ:��p��s��-ݻ�:�-�q���4���d��^rL �:Σ�:��<������s�F��׭Ļ;Ⱦ�{Y?k��0�\�rC��1�&ӄ �@�.�<=?742�?�x�j�_�f�^� �Ex=�8�EO`�-���e�W�2�Qm�Y�x����@��633Ǔ�!���,�|B��!���N	jgQZ�AV��<����y��P(Sj�M�9���ůwSl$҅_Jޭ��~S]�ϫ�gd��O2w\��wv�\���X�W��4B;�M�ԝ���yǳ�F��{��{�����VR����
�XEmjｪhk���,j��ڢ��o�v�Mm��y~��?��_�}]�|���>׹�	��%�{�O#Ϻ.ϵ�V�Ҹ��oNVݽڒ����Ӌ�U���j�
���$�J^&}y9���ҲXgq��o]n�D��E��O�l����W��D�8%�~xV�M�����1�!�G�ز��h���7��B���#��^�V��fYM-���1�C�$�m�سV����)�xN2}��N�����]e������䙓�/[�IN�����}� ��x�R��:���F�6C�|���0+�<Ƹ�.��>��	R�l��%h�ݣG��{��x�I�ektO|�}i�|�ko(����y��Fs�&����NQ	-�:���Wr������g�	Z�v��P�>�_e7��P�`�oX�m���h�ɒ���3㠮�O�o��E��I;����w��ԝ��I��-Ѝ_��%*h.��c*��x�ZRy�M���c���7aץ_�_pb��Ϝ�ihh��#�mS�K^��!!� /��!�%�Y'
�v�U��7�>�v��1�{��K��D��R���El?��.�f��}�H��S�aB�E���Q���!g*8a{+����v�v_D��\CsH[���c�pbK?��tz`gL��qvp����1�׶��RDcc���B���wG��yhD���Ez�v�1�ޭ�.J�ޭ�p��d4 �cvw�*���(lxiqQ,|g��_>4�)�A���\������3�$bݓR_�p����o/��'lE�/"���/ƶ.���K:U�"O��{�S��1�y����<}��ƱN�Rlo��=�#ojR&��O9�Ύ��=���ˋǝ��������S�׼���w��.M��d��Md�?�s��������zӈ0����ȇ,++�8='e8e���6��ŕ�b'�E3�@t�9����6*
�J8[������ǫ���A�ю,nP�T������ �Q�m�Ukn��瀎��5�f�~u�2?)L��s�0�Xq�A��m��9Y���;��e�Nv�X�x��\D�������˹����79o��{��4y���8��?г�� ��8L��`8��&�tE�Y��&�Ϋ>Kg�y�C�	���o2�4:��0;�Mvʸ��ԣ<��p8����x"0�^U��kO#�
�W�i�֟6��O�.� ���ۘA�b*%`�V$�M�}�y��,���8��0�̽��k�����-�H����ጪ���dzٍ��4q��)����D���,�7&c*p������z��f9���g:ތvh��Y�ʩ�n��Β{����U�!eb���Բ�:�U�pn�ϩO�'c�(3״PL�JJFI��.�������p�����~�����<�{WVqZ�����B���vK���'��n�hr���o���_4�3�t�˖]���YH�>���MMחqљ�W����������,�*�'������k�y���.!����kꂂ<�4����Z%�_8���γU9~����v
&#Vc��7J�tɏk>��4�Z�@m\[�qnUNV*Ys/�#�:����T3X���r����7�q�,1Qo V�9���mv)��Xoy�x�ƃ�dOMGɚH��rw���g_����h�Ǐ��%�\�4<vID�W�>����Ni�w���/2}#�����^_/s74�N�C�������?6����:"���sx�c����Z?V1��7r)�xR�x���U4����gkKn�|��,p��@@v�_{��t*�PĖ~�ã���~<���[ۻw�������oA��b
�o�B�D~q)��ھ��=�NI��u�$(��)a7��G����_��f�]
�q�ˏV@D�4�AZ(�xPry\�`�7��\��싺Gs�� /3��/�ϲ��]�|��|�DP%%�޿��7}br��ֶ{4@�6�5�N�r^~��8��Ϲ��Ta�9Sx��wFF�,[b��/�r��w�y��Š��=���5<*Uj��pxZ�-#����(�.���fO߳*�wF�si�X�L݂��'�J����S�{e���0*��-bY� �?�J�.��gg�p
�9�;l�#�p��X�I��86v'8m�}v8?�ئ,������!��>��l�~z`rRLe�?�S�����_赃R���<ӫWň�̙6s���$yI�s2�]y}����ݾvFf|*�1����(����	��27�"l��`5�(�����&�S0����%Be��(	~�r�O Á3�	��)+	j���AJ/u���c���w�b{�+Q=������Q�r����Q��<�b1�՟�V^��3��M���2
�v�����t�h�;�(���fp����k�7���|R�Q6c�¼���5���E 	W�q�0$@3����5��/6[.��R.�#4����k�;Q �$_H��c�f����W��t����(	�E�?_
8�"mlpB���	e����@z	AA�`�l�?{j{�s���2G񇆺}�MF=���������%b �M�%f��J��D{z�_�oo��0�$Nq�8���UF�=EsT�[O�`�+O��a��(�F�$���be�+���Z�^<�V�%�5�(-s�w��2�����J����B̙�$ӽAN*��
�dN�'O�>14��p�Ř�ദ�إd���܍P}��zy�e�oHө��PjB��gƎ���%ćN��fN���dGz��~Zh��CV�o��$���lI�����Nmn���;
��*�ܷ�!���Rg�ۼ���{�wsv���1hFn�"���XC8���pH/�KW�_0��hۭ$�WDX�c�3g� 0bÃ�1"#�Y#.�*&���F :I��L�h3�;(K?���(�?�������=x�h�hŐG3����z���t	��A�
�t�"�n?�e��H���,+���5 �A# �0k��s��7aw@|�T��9҈�R�D�1�X
+;-�!$���1�j�7��l�S
��@1��������.�W����D�/Uw{���"b�S� ղ�<�D݀@S���R�W^�$�� 8�ҝ~{F~�,Mն��\hֵj�>�G�#ωB��m�CCh����8����mP\Y��<�3����:���a�[�y&�$�j���m�t�imH$���׍򗲐��������I!�܃)i����7t@�VD���8��C0E���W5N{_��7��=`8%-[[�>w�ƈ_|�Y�F�.~<1%��3m�$�guV[��>�Wن%��M�_�8��z9�e�+�4�����T��Q
��䎡�r	��TX����!?�;�QuP���R�;6�"@�W�ajd�O
�
�L�C��|&}������/����4G��l�vPT�r�qM�&?k�'��S���je���t-'��n'V���"��h���hq�sI >�䳛��4��{�c�~`{4rxU�ǁ�zqRw�G���r�3�aB��,�v��Z������7e�x�{\�{��4��e��]�_�� L��*I�}p�,n��_>0A{ӄӡ��?V��HId��3O�(<�e�A�V��M�q�<$��FF�,UV��no�' ��k��ɣ��i�2>�a�H�z+?KR�Wt���f0�S���nm]�t";*��������ӧ�A���ǻdo�xɳ۱������>=��Aoȥ2��?�8|����`}� 3���r5(/%t�٩6+�]eS�zU�9�Lx���5�df@^��*�����\6�ؠak���5V�u�2?z�AGQ�@S�0��}:^�K��uX-#�����)D�D{��-�������Kg�h&8������e�Oj�����ӽ�����0�u۪�}|���z�w��G��H߈��yVMn�%��c��$�o�v��,0śJ��Lf�<�
l�r%l�-���쁌�u�l��T��NLy'�E>�WA�SGB�yj�˳33�qX�"��fYqT����_��a��^��e槂Jۧ�|`Bcj�o�����N_�+5�?ݰ�����"us����[D��cߺ%� �-J:N�*b"�����~8�:�<k��ޟ
�Y�g�&���cP����R�q��=���L0
��<}��E�N�a)o�S�����k��M~�TFg�?;չ��#NW)��\��rtm�`�ݿ"S���f3����Թ'�/p|�����$����W~�U��R��6��Q�-=�9����aK�r3���v.Zi%����ʋ�~R��2t�x�����[��)*ll��=��.���j�PT$E�w���@���r.b`��=��4�"M���z��RΆk9ۧX�:7��}�,�}א3��7B��_���μ�z�Mi���S�7Ҍ�̫��V����F�ZߛY�ٮ=���OUK���n�#�:*��m�E#��ţ���z������ Fر�f�n��\����=C��sbӣ��Z%�Au-�?g�Y�2dS��?�N��k��	�8�[�r�	�}4?7�4t�n��T����ş'$AM��n}����ڴ����{\�z�x�'uA�L9�2A��l~MϏ�3Ew|�=?b}~0N�P���a�w���ݕ�;�xi���8�[AAHdX�$K\&#3sVU�bj$2�ǁ��8\s{���v��~��@�y�´�B�U3|���trs���khY3g����}���uD���o��`z���>h�`���<b��VY�'ogM�B1�`H*���}�#
�}p�y��x`����67^+��$gcl�*zU3���d�d�l��'�q�&��_�t������x���a�x�'w2�h�m����S@L�;��)�|�F(��ձ����L*��L��v@�୏A$��`��A?~�쉼�7^�8뺔��֖��X9kXlJ���4(��������&��ʝh"��?��pԚZ?rp�	n�H g��H�^I����߿���](�t�{��S�J�;+��~���1i����R�~�<(c~�ƫ=�{y�CD|���Q��I���EJO�����r7bD���aP���
8�1���6p�2�g��p��y9�v�]��w����'cX�z,���=ۊe��g@=�C^��L��@ꠤ�n�o!�N˧½/>_{0�󱫽��1}�2s)��y	��=��Ҵh�P6�]�<�j����ՙ8G�{<?�?;���� 8�O:h�����6��< ����̃��_�T�o㐠 �(�_�=�,�L��u���vRm�鏈Ź|���;�kǾ� ����s(�FVHS�섟%Lz��Z|�tKC����:C��9DPZڎ��2Fb%��[b���k�S�]Vq=�� �v�1���M���A�bq�@��{aƶ��8q3@l�u1,��!��{{����Y�2],��8��k|n����}욯h�x���Ǵ�(�}9��Kq�O�����q�TU��vTQ[WW�xJ7-9P�]��S-� )��'Ѭ�z�+2ǲZ{��J��C���⨜蓼:����-$#1�a���*�΀��.p����PˉA7��S @9|�T�������l 1���|Qb�L��5�`C�Ā}=81��U��i*��g�}�N�NN��h�cj��'^�:�W�T���X��~<���0�!��!�L3_�������T�Ǚ����q9F�_�w-�e�n���+��dK��=:on{���o�z�G���ïְ?M�p+5��J��(����ԏ�zh���}��I�o�x�s���X�Ć4���(Fة�Ƈ�L�R����y=�ɤ6��0
jts	�u�U3rl7j$~ɪ4����!'�����ܸ�ܡ;�s�,����Z��j�Sպ�?6�@�/"���y�=�h�[�UN�O�����qY9v�|p�9��_�'�
������cA�q؞�l�6%�<h��X
U*��pxs�xv���Y�E4�8@JGym�����h��N6b@֒� ������x���+�������K���̲j�ߑ��� j{�0#����e��WJ��g���ɰ���È����#]{����s+�v��ٱ1WdJ�����(�@·MԮ�P��]��#�lv�� a���c�V�3����?�h���ȋ4[w�[L:[>\{ܩ� W2�Uc8�����&S�I.�[���:z�����x�ߣ�u������t:2�uXi�5`���V�����F�1"܁Է6)��$z��bNq����ؔS��-Ǹ�4d���j��]��@�!�@�D�c����D`_~��ɉ��+B����� ��Y����3XH��Ӵm���w��Kd$�c�$��|���p�����0Bh���D���N����y�&އ'7��ڄ�����&�вs2�§�!�!h}���e�V���9����d�&��ϗj���P���C�^(L����l�Bܼ6K�U?�jC�����2��}R��]gnP��
�g���:���5ˉkcɍ�(�x��E�Ҽ*��lɗ�$	���\5�M���B���T3q�4}��|�V�$��:<Y|�"�۰%�0bm8� f0�7# m�}�:j�~�1Kkh5���v��hTڌ}{��+���#���Oob���x�K�i7������Cgh���$5׃S������,�l�YH�q��q�����[F�~qy��������.�����UR��\����LK�2o��C4� E;Y>���ד��-�P|�o�x_:��,��zj��,ZP�Mu����\֑���ڔ"��>>��zw�ܴt�+YF� x�K���i(3�����*jʕ����7ߚ��7Sc߽9L��䲕<��A����X��Uz�D?ak�utt{��[%~���h5�����FA�me�е�3�T�@^�mM�ޤ�������+hĈb�����M� vqZӜR�������_bF�\^z_N�m��ڳ%h��^��3畒��Na������7<��<�*���~�Ʒt�'&&�/�P�!�[5w9��j<�Қr�Rt/�<�3��	�g6��.�-�2��u��q��
ׄ��#��rM�`�!N��Ƙ�T��>Z!@T����r�2���w(xʵdm��r'�A	X���1Z,�
�2����T�T�a0�Nt�jcP)��ț�ة&v�VR��N�5ܐ	~�m�0���5��JM��~("y��{�F�S�g�<��9@.�ݳ�eXق��<�)Lc܍��7��>m���U
�F�Sq3s��S�!�x/��m)M3̱yx6�1>v>��`q����b��4��G'�!�l �b�
m�r��x2tn��u�����q*Z��?����W�J���}����	��e�9y�V����ͮF"ErЕ��:g�A��5��Q�,��*t��[�Ȃʲ/�󌷒��
N��o��[Tڌ��'}!f0�mx�4��{�]ا��i/��U.��)4�P
��l�W��^}��U���TY��x'Aps��i��K�`��B�f-]��}/#<�T�g�&?-���[���)�e_�٧������J�U^�J�=�n�|\k��h+������6���"����y�D.����S^ I�p_~ �������Z-2�c�Ql'��lZ�R�?]c������gV�:]�)�&��S���,՟<u��"E��w�W����ŏ�	}|�G%���XXQt"��8G��9���e����:ȋ�}����R�Xŋڐ�7�7��=L�e5%�=b`��ો�M�C�3U�hH>�w��NA�t�:��2uC�%��E��$�f�=��<7�P�豓Ra�ϵ[Y$v5b+�&6bJ�_������<�9$I$'S�j����H��e�"��]G�v�&5�n��x4�߹����ղ�$�
�9�����FVzFÚ�S�>߸�4A�������#�M�3�ɰ�������o	WV�����C OV��	�oB���P�*��}��he�K+�s�j��Fp����РPC�h��m��j/�9��N�C��X9�n}��1�H@9��vV�T9rk���bd777��L���ٟČ"�\�9_o�na�S�Fv/��7~��(��8�/�C0�lj��E��/v<�U����}� ����1/|�=ݓƘ�lm�W} ���X΢J�~��[����=�O��(T��j��g�P�#r`��X�F��,�<Z,��?�nVsod����b)(Z=7ߠ�b�6��ezuĘ����� ���K��Z^o[SF�ލ�u���8�����/� ^ ��sX����S8=I��� �>�jV}�~&�ɝ��6��`��+_�`PX*�����S�LkO�nldLA���R���v����G�K��9q����Q��.E1�F�>�
dh�ewT�"2|�B��R��(=i|=�sO�N��٨d&��6�ߓ��د���$
4o��	��=P��f�4�=�$��$�d����ٛI �|��uf�/��ȣ����%0��MPPpy�Prr���[�'�Ü�E�f�y2o-Ϫ&#H<vD��}��� {g��7܈�oh��a��r������Ō1I��G>Q����=,'�;�_������n�d�� x�g�_�:5��I��}`Plzt��ׂ��齅-[��8[�
z��iF�v�#T�{�2�7?,��"x=GX� ܾՑ���Fl%�ŋ�7h/���d͙�_*q��P��s| �u�W���(z�>92���-e�t�\��{�H�R^����9&gh�7Q$��sh��8g���ޖ�Y������n�6c��^���M�K�Vuyì/���ҽ̕����j����$ml�e���ͷ��9�&pleN�ڃԐ^K8��]�$د��ӅJ�6�	�DcC^�|��L��Ja9�J7,�+8%K���Ӄ�I1��>�/�8Z���f�C�,!��Y&�����[9��f6p+�M��Y����hs4�L`�U=s��0Wݍ�),&�I8�����B�Ĝf�$����o�^0s��J���g#�`0eN>ɝ�˚e!��nZ���>�}`����Җ��uQ
��W��G�A� >���~�7ߋ�-Q �_�2]
�Vo�|�����B9r�O�BPq	�Į�׌��#���J�Xr�EF;�vC͏:-Ft���e��
���7ҷn�Kt��a���A��e}���¥߿=���a>�I��rӆI�a��E�〇�\q]{B�����ׁ6cn�<d�eI�I���hZ�N7ͻ�O���2&��`�n�7��O(Sр���X�:=&ѴL�+]#c���2���HfZ��O :���Qs��J�9FL=�� ~�����'-��52�U��
�4��R��p@����0����",���t{�HJ)g�;V<�[ ��P1��_/��߼����+F������s΍�p��:�P�g���Ǯ|��b�����<���Q���°��R �%c~.[�E=��)Q���O@�v'����Ƅ�/��19VΎʎ�EV1F��m6Wץ�-�
T�d8�w����ӯ�5��x�E^��f�$�Q�@#zlY�Z����ő���gK�^�ő�5��RR*��V`^EV7Le���|����O�ʴh�O�[�����߇(����V�j�di��k2�V�#@O[�`h�w���_/�D�5���o9}�MEU��S����嘫�T&�2 �1�<d�ksß��W�6��i�[��s|�����Q��(q����"�t�ttAq��\�f27���{q�ol:���,Kugw?���z���5ْ�`B��a[�%��Fqt͐�Ov���))0�h��u��.�4g��(���c���C>#�dQ֌S���Ƅ(�����q��R�-UT����	Q�3�|rf� @�V5��8��g�^��M���P�y'����V H4*Kj�s�Ĕ����+�T3��9�Z����F�/�1��S.�����mv)��)��u��5uK�+0��x~��f:�`��_e�p�/?#�8F2/5��R�E �	��F&kkdW1��c�?=_�aХ���@ӯOlU�&D�-�9qPSv:L#�5����Ѳ��-���'�1)I�66�dQ�pr�<�ttW#SPY3˖h����34՛���Y��i��?t{շǊ���l��ٶ����A�>�U���ҰV�cé�hq��2��\�=���Ѭ��)ҷ( ��O�Zj���2iY�?;AS����m�e�Қz���+W �Q�W��1����|QtԼH�� �����2�4c-��ty�^��=�)С��<¨�i�X������$~G"ЀٖC�L�Y_�x�n4`0�&���r�`)gcQ�:��JeE��P����i}y+�[Qn���܊RT�,U�B�ǽ5�B~�)6���G��vbL���{ɒ`��*��� ���4�T�,���bzi��ϝNMr
<LrT�B�>I� (n��䩰���\
�5� ²O�s��.g�W� �BQ0�'  ^cx��G&�!Y�"(u��}Ǖ�<I��ڡF�mE��h����6/Z�7����M�b�N_23 |w�6O�A�������T�utX��w�=>y�Q]#(%N[�W���π��-}�����n�+�++eՌ��y��C��SS��]�*k/�V/�m����h�j�_bOw�3�iٝ2��a��p��ϰh���������/R��_n)]/�(��P��y���v��o^�l��l�'��+��G��a]�#1
4������y��ک���a��dAB�Ĩ������M!���>s0�hxE��r,���%u����]��v'�̪�^��`+�V�?=�����`�j�L��;6D-�Ll�n��H<`Bo*����&3Bw�zF�w��>��}hP�J�'�:�t���.�s��r��[����j}�ec�F銞p�)�@�h��ܑ��&`n�J��	�?���ʘ�Ȃ���j
�و]3��XK&3r���RZ�W�d�'q�����DYSf=��Ov��
l���7UNZ�e��_<���/&�1��.�����^�j�PV��:\�Z��O�o��,���r��d��h@�����say#����U�'6�`F�}gcb�Y"���|�B��^x�"_�̩Vc���,E>sSc��̦����Etl��#��O@Y��:��o��Z��d���Ut��0/�9�%K ����݊20��^����	�tϲ��O*�n_&=+��O�m��CJQ�.M��˰k�����I�q���b����	�?9����܊���X�]���S��?I2
�*��c	���Y�;ΦXU� 0o�{<8���Z��^�,����܋��OH��_����nE	R���
t25�2^&|sRc�3�(�V�Ùy����=����.�8:S�qi.�gM���;o���fC��%%�>�u��z诙��Khbo�"�N�]{��{�Ѿ���xxs��x���ڃ��\��)
/ν�Ma2���ˡx�)rÃ��v
+h'��QZfD�1�%�՘��~����|c]B��պ VHa��1�W��;�Jʈ�E���}�g_n�.�9@�Gi!�w��V��ӹc�};Zx���� Im�����$&���j�c�����A>%�b����~�Ml��r�Q�����jd�/{q�W�_�2^1J@� 8%����}
U�v�Y+�p�_�>:�Kq���MS��Mcg)p�?����,B�6�~���M�85}G
�CT���U�/@�"H�u��}M2Z4؀GUX�C)C���uf�@�y§�y���#~�;���)1��j�&P� ���U'����C��N�c:�g���)9?Ʊi��m`��M��	l�N�F]��������ʶ�P%
��n���s��/qQt,z�`uj^�j��ts*���R�u�>/O?��(W�O��ȼgZ��V�G=��jFh'�p��U�^��!��ܹogU[dw)8���5c�:ӄ�_�[:R��9�68���-�2xM�Pd��}"���gЊ���þ���6v�{�[-�����+��[������X��25�ύm�x@��;,�D����vfCV�7T�NY}9�4
� ̮�t�3�9�XV�������
�?�.[�����O4�7[���*
N���ع����+7g|�Ҩ�� uu8
����4?��K��j���o�ݾtZ�a�TzG��e^�|��-����5�i�-�����1�8Ő�K�����i��k�!��Wh���R[�|}}˰�9b��9�1����`���%���o�'k�K�/0�����E�
���o:��`(���9� {�����o"�'�}A����gbd�wN���T�b0_A�eg�\k���u��
����JUInc��
����fBT�T�����r�7s��[���T�ܺ�ؚ�����+��\�[�6��I*�C��wW��n�Y�g�w�*_��{B18u����P�����5�j��Ó�=��5���P�5|������ؐ���K��ϟ���"�I�W<'�[����v��{"B	Q�^�v0��뚿���[����Ǿ��:�P��3 �ı[����i\�	L�#�H�������vR�MC�u�'B��#Fʍ��69H�����8��z���gB8����M̏�V�y��Q2�����^�Z?��nJ eJQ�<=�1>��0H��9M����JcĐ�b�O���de)fz�;v�x�[���|�`8�W�c�wF���Z�2Y�> �G̩U.t�{�і����v^�g$Ro�����Q�J`#� ʨ�� =2��(|i�q+��ڨ�ggp�]����0D�4�
�ƈ`w �u�y�>$q}�aN�G�^g�.�� �]�����U۬ȟ>�Vydx�xf=cdU�  J�ېZT����R\/v�(d��<U�����_*�? �Em�}��J��U����@���؋N7����MH�P����p����?�*���g���Z?�
�AY�ju�"���a�T-0*�Ɋ��W�(��f�c��)�˟�O}a��m��� ����	�ʡ�*��c�e��^���ڀ�;|����Lc�J.D�S���<�q��v*�b��Bd��f�Z�*�bu��b�l���=T7�9�N޵�y��A�����&[X� k�grҦ�>�ȍrd�qJ��퉲�GX4��;�mO֐sxuܳ���~(�7���f}t��A�bF�9���sҟ9���7N$@x	�ao���XC��yȇ����RC)$3��|m�F���z��6�X��ʻ���~-���������6,_khg�Q�fг0���u���R�3o��+��$$���^��� �J�>���2
��*�ڬ��-�'2�B^g̪��ݒ�����Ɗ�7k��1��zݼ}�K�9<�.Cr��j��2�D��(����gU�L��.�o�{��T��>�ia�����<�=C|���� Jl�������
K6j�>5���*+ێ5�_,MMֺ�H���Y�>pAY���θնu9�@�}��LJls�w;k�����aZ�^�4�+7��ƽ�z�Sׄ��<s*���Ꭽ$�Rx��`O O�NMeZ�P{~`_.k��eOڱ)R�*\�l����ʰ�r	s�X%<|���2��jN�~�����BZ�k�"�µ�7$�I-Vk��3��U� �	b�D &��b��c��~˼��.a�"�	��+�9��'�b� ��Ж� ]L����K�*�R?��Gy�Ň6�8@��b{+����7�P�O��^=s�}���Ljm��_���:��;=ʇ<�����Sޥk@�;��)��c�������k�2��Y'��|��c�^���ڤЉE�Lxi �}"��v��iJ"N�̩�BP�����q��x��E�zˤbI]��٣o�#��J�]8�S=��*�#�=�N8�c ��i��MA��)��؈��Ń������[�|m��~!M*�aV7XF�&6Z����aVϹ��QK��=ص�W�K�i:�G��^>��%X
����=�O��	�\/F>�ک.�7��$�qk��.Jә�Y���>>ܚvj%�^�cv�akd�1e���A��sCP�A&��Z���]��ʕz��R�v�˞�������H츌�5�z�a��r�k�ao<��2S�S�?�/+�=��u^�
�%,,|��9}��;�_ֵ�yY�u��dX1�[����m����x�p��jd�SԄ��V�X�SY�0�2�?{j�k|�n��]��եb�Д��TGI1�j-S}�p��.�A�9�Y���ʮ�[�@�{v���:$�T���gF�O���ﻼ�zy/�L�Oe�kLإ�����؂ (X�m�u�t��3!�ybi֥dT�����7�zM�;8�F~	lE9���v��MsDa\o�p�tUB�{��)i����y?��~�`�v*��v:��(ڹ�q�Я��Q�%M	��/9��K(~�R����'a��o/�������}�G�]F�#��=TGFi�kFl�|���$���u*��JH��d�dɦ�6C�'��@�[���j�i �S���e��� 8��)��}��F�Z�(T`��n:���T�*�)�^�����c�O��Xt*�N�E�[ ��{Na�r��ZUe���;�q=��aHR����Q���wJ၅ {�����ڥz�������L�vƅ��G�ٴ�RR����Q��y���O�D~ҧ`�O7���ݒ��ͰH[��+J+V��l���V�e�H�U��+���}�Z�{�+ptt9�|]hT-�M��lY�>G%e�s��=P�}ho��9�O���:�?����E�BI-�^��.e+յ|!��>�5=�^��u�+_�Rc|�������ݵ2�@z�N�E��w�,?�An�&�
0�=������1����b�s+�����9V��$ސi�����b�{�Ԝg YJm���,ΐ��-�|��,��-���?:K����U1��&�4�3�s�(݊�E?�AL���
$<�u���W#p&%p@�c{��"mK���X��2
�_a?ݟ�7�2�}d�(;V��n��<�P�wh'U����	�؍-r�������IG��Ȼ���/[]�>���眣�C�2'ax˿ RC�k�nZ�Y�p�|m!��i�-�ϔ�BV�
�w9�V��S��\�V��z_���v�xڀ����}-�<鵙�d����0L�k m�˂`xaE�ꇹaCk�#U��ä
�` �'�~���(�ADh���s�d������k�=������a��L���WΦ�,45��I�#U"�lQK �S�}�B*LTW�m�Σ�?�Q�q�v�ǚ�t�y����۰��ѳ����c�_�m��ɥ�xXm�����B]��(6}(scY>�Hu:���S��y1:z�wkc�� 8����y�Ӊ<�|��LC�w@�S��H9��c�q����&;`<��Y�˹]E�y�\V\7�*��ӷ��2ʢ�����a�� >>�H����hV����c�M��O*��/���$��]�3��J���Ɩ�)8�H.����B�&M�H�nG9�w:kk+��WJ�[&��)r70CS��L9	�����8(tg�����']�3�n7o5�~��-v�*������n�ɂ֫6�nu'����,�jʃ�2��5�ۉ��.�,�x�-d�i*	2�i��b�a�z3��|'��}��*��������7�g��wR��{��nW�Ӗ's�&׍��R��oY�����ݮ�����(-�����:�c�+�ԁ�`h���qt�6�&�ż���Ƭ�3�7��G�k�؈�C���� ��A�0�DfD=$!Ъ�Bl�8<�g�m 	
_���L���f��d�Ku=��O�(���l��;dM�R�hvު�s��'?�q��ߓVS�:V���^��D)�|j/ޚ�����4^�2P�!l>kwHP��?�����rT&OEԥ���l��Bc��M�U)Ҍ�(�S[��DGa�P���E׳��TM�a	������S^�$1��%ܨ���>X�Εi"�8�p<൨3�~Zq����S�Ȉ����`fB�����]t�&���hS����*�m�t�y�!܎��r4j��SשWK��0<{��}���5���P¨d8Q�0L����q�E&�âr$���Pt!1� ��f��֐��� j���u�C�[��I��a��
�	�V����5uVh����%G�%=A7����:?n4{���Ɗ�>i=�*?�I���xr��|�>�s�`�'�����&�Ճ��~��Yd�6{p� ]׃�]�����>��pYs����5MX��������{d�4��5^��^��a�l���F��(��o�8^��#�6�i�<���ߝh��i���jnp��ֽ{�JJ��>5>�*4�vH!;�?,]uX��ߥ�K�э���0��RC�;�S�ѣt�8dH�Fʁ#DZJ$I_����׮���9���|zP��)��=!qщ���_^��}�����t��f�K^V5&S9�B�����^����I��zNۜQ��7�%�"f��Gꧏ��b�8u(�"k�b'r�$�W��GKs�}t��0iN.饡��1C'�1T�a��`�.*&�^J�& �:G�8�z�뢚,���7�W����%Xh0Z�-͓�~^�3rB� "��u�ju�����+Bq��!*��ESS*�*�ҙ5��A�e7`���a:n�_��pų��x�G�0��գ�}��WU?����<���x鑾;�����b���`˹�qx�d�f5M��9�XÐ��pȇ> �Я��-�\���\���H��I@�1C_������_��#��[3����'�� �캤$�+��$�Ű�]3�rPL���0���i���fc�M�~V�`V-,um���Qĳ�F��q~��?m���^��P:~�U- ���������!A�i(�a���Xk�+	 �x�o�罖1�<�E��7�����P�hZq�
/��sJ���v��N�<�G�l��\T��^�4,z[�'EĊEy�}f���.��sޡ1";�M�sC�ҫ{��J� ��W�񀍞��?f��ɪH�dh��;�j�g>R� �ب3�R��=��8���^��۽ �_�;x�%O<>��9ʏ"��d�j��[�]ۿ�_J��~��I�p�{+�JĹ�g�8��c ��&з�D<�Ոo�+�S�X�X�6�������%��᎙���-5Ն��3�~	Spn��lܯğF��r30�Y�
���߾�f�5¦�Be\A��|�B�Lq$ XzP��wJ.\Ь����3��������F�	��m�bA~�{šq��7m�zD��7Q4�y[�Ž�KS6����e.S�"�q���:��o��ڏ�_�c�b_;
�4�^���KK�8�6�T �N��G���9L~*^���3�2���$/�!)�D��U�F&��fs8R���e�)k:-���:�bXP��Eb,.�o��6JM�C���?1�:��L�~�KS��p��)��sL���㣗=S��.��r�&6���oU�K|�4���Vsަ5�ː%�_�����*����u��u��byT��~����]I�w�u`b�g��&���l?ό58�ꡫ�ņS���s&�M�����l�Bm����Bܦ'b����lG���L�<*���� �Q�#E�%�~�1��)�B������7�x`p���c�������b/����w�t�V��T[�BK�O�����?Se���jh �����v��|H���y�$���:�0^�~?���{��)�1(�����4��z��hb���M��#�>R<��,U+�j��2e��
반0�s����e��u��`�{\��s&X�M����<N~�J+��N�G=��-;ö��|�޷�S�J��)�ouDz-j8���x�5��� ��r�$�վs�Vʪ�4l@�b唆?w�_0+CWZ*�Z2�=�|y4��eDR^�a=L	@�`
QTT}�ѳ���2�����h�t�g+8���!�d����ڌ؟�h'{�i-j^���ڑ�$�N,S��a����G�׺3edP�X��:1<`�:�#�{��)�'2ȓ�r9w�p��\ٹ���Tv4?mѕ��N��>�~]����� ��Z#���,���o�J�5rvi6�/�o�!7�
����}ms�Z�p�Y8���->���$A'@��C���͔m\�{>_����;��5��l�+G�=�n�D^7�-�|�9��h�;"}W�j��?��\����ĭ-�A�<qҼ���j��o��J��9��%�JT䟦;bY��Dt���yp6�������T�t_��׳��@J�"���59�sxC���Q�qPꮣ&�8��CE;�]�08��U�QD�cP��q<�Õ��5���Rl���>�F:�m�ˋ��ϫ�3�&��h�����ٌd�
�x���I7X��%�}�섮�YC�mh��̈�ef�P�H�|""� X�bW���Z�P+���H�*裭�\�8���6Jݟ����I����N���>�$y�)�3{�����:�]�!ض�A+�v?j�����¤���C���qy
  .�^rUV�)E�Ux�>(@��Ub�U�	 �`\�{�;����!eȃfV�"*��Q�/��8�á�S�שC�ק����=�+��K/�>�a���(��8�E��n��Ⴗ+���?r�"�����UX[t��S<1�R6�n�U)`���n��S�{C���0��?�:5�7IT�3Ը�_a_4�3�]��Z;HvL��t<�}�Ɛh�1K��p�c���M�ʯf,�$x���Gi�)��V�Y���s:�[i��n���*�;���hP���o_���>3Aw72��ׁ&��٧;rxS%e��?�m�������+�������}o͕�����G��e)���.���cɄ,��B����GE-(sa������?�u,z �'.z�>.z�ʔ�3�$�F��$Q��Q�D���ϿV:?������*C�
�]U�ew�<�.�6Fb]ެy����;��0gMz��ޝ�zW"����ڗ �7?��h3��Ҡ������gꄓ���2$h��Z��=^��*��5�jd.q�+�_���MD�lh{�$�9��U��B�G1��RѾ��B�@u�h�<�Х�7�S-˞�-+���0<�jK̔:R�9fF]�^H��)ě�T8H37�5�	��c�se�Oe��zi,�*<Y��8vX7b�LIDx����K�!l�ş�f�g�ޞ���n�0�3"�O#Ef�4�X�]@\�=���	��h���F=O�A{��egR����ֶ-������:%!We!"��i(��X���.��j��e����5�Y�O�M��H9k{ڏ��% &�k4�*ƨ&	w��ڂ,e�����^Iuޮ�wU������;���h�F��-��i��ü=?����֒��dZ��#	��7��r����Rk}g��9�&ω�E�a�����u�/'�_ 0l��걸��-6Mvr�aa�0������_���y�[�2��
Qu��g�ϝH��8���$�4:.��xk�N���?��^�����i���_��T�<�[qb�q1nX��}X�;T�0��!�J���[�<q��ޅ�|q�%<~��n'<��rBM!ʣᶴ6PPX��͡&䍉�3�>z���%Z<��4�i��Ij��pxAF�M��>��w�ӗ�dn3�?�+���e�+��=���k�U��:bWlan(F�j1����N�p��}����G����)\8��Ս�۾��]Y{f*����#�K^����,84�&�%���JJ�a��(�t�*�g+E��Y����]/�Q�ȏc�T�7��ԉ����1�&���5p�����[_��/���ԙ��R];p����wq��Cݜa��;xb���.S����t@��b �MwP<H�u�B��Y%�?������Â2Ԛ>�>��� ��5�h�&t��@���M�e����:��b�{����$;�ΌcA:��wW�è�3���M�%�2ɾ��bА���X.EQ��f��G�PR����5-OI��}aR%�Y��:3(HiUm�B[�%a�D���?��g�f�I�"2���z\�;$NS��,���a���0y�_\zц)�\�
���t7��H'��W� D-C�ʈ���-=���  H���d�6"�^1�Z�uz̹D���=�ٮ{pӇ] ���9�����SY�����o|~lT�>��0�2� G�~�D�)N�EI�1*b:�Qr^ǿ��G�Q����zB��j�Ks����K�ݰ�]1,ݵE���}���D�Fw?_e�/6�-���}Sə�e���5�%����M���ξ��#X9C+�Mq��:w��^�ȳ�/իrP�1�Ƿ��βt��셥���e��#���Y�0N��ɕF�85�/O|W���%/K�)Զ@�:;7��3Qe*��}8�*W+a&r��@J+vҁ�}�g�Z��1�`QMt-l��k�zA�����s7���2;�Q�����N�cDǤ5!�.�DP���L3�3A�����$t>}�g^���>V�}5^�e��l#�}̅.���m_��w��35R��N�tp�Y��Q,B����lOL9�wŶ�����]E�(A�(�i����%����h���:�<�$���տѝnwĉ����R���r�6�>zFB�xn!,�!T+*�շ2��y��Qi��h$�� ��{�-]�%��Ar�*�IgӾ����l]����MbbhL�󃴆1�>d��E���k"H%`��x���)?�<a|��X���\�k�ߠ�>�l���7DS���'�~�猪/��슞��Ȭ�E)������#ڦ>/�״�E��A��9���vVR~��퐣�C�/B�5�k#B/XnZ%0�I[���V�|B�slq�#��6s���=i2�8T%�������B�JCԬO��������l �]?Kt��4�I��h��;����mdx(�C���<��E���,�������-�M�2rԦT2������;������c�l����BJ"E$�7���H���Cp�|�V�J����5䣯&�D�8��(N�?^��+ r>e�σV�۷���w,�]��5c������iW�799���*������Ҳ�L�����&G�B�K���It�fē�:�.��r��>��U�A�FR��&�vK�:ƦNM�����\�󠠰8��8tĔ�o�Т?ġ��}�r�P�o�EV7��Nu%')�%&8�-�1�����ҁ�i���:������⢨PaⲈsA�������ڈW�����"��s�E�Y )�08��-Wt\��%m�d��Ոo���u}�e������
��ۈ�뎯y�@���v��}���oo�$����E�#��E���ky==�w����G*�����<�"�/�tN��f�?'���1B�u������ܝv��\<�0�����n\�lBI���|Ss6m��>�ĳj�d{��'�]�r]sE����oNBA�f��ר�ț�/9��ljP��''� TީԿz&��nCg�cOO}��Y��H �=K�#�=�k}>&Q���Z�zB�D_�Wy�sxi]O��b��i���Q3�LL:� �m'_(�w���c�����cTV���i����Z9�@"��$f�5��l������kó��(D������6Ӣ)����U-	1C��żr	`������=EpA��v$��*���Nn5������5m�\�[�yER����'����KH�\���5�*����x���S���+Sz�$5������#@������� �s��K��Q}��o]���G�ԧ�*;U�0�{�DC�sE�y@Y�L��"Η��� �j�=4g�
Gx�1��s��ւh�`�3�p��3�� O�t:iČ�K�
�}j�;���+8�>۱4��vQg�2?3����S��r&���h���t���
���0k�;���`�(h�pfHs!H�@�i��cY�&��F���ZƎAA��=�k�)��0�Lp�V�O�FfYi�b�v25�/*ki�*�x?�B�� ��&yP��X���Y_+��򧌀Y�:(yEe�LW����2��Oؾ��Bq)��.G�1h1�O� ��ggq����q�!]�;��j�!Zy�Yq�8縯�7�/۾��� 'y��x��,p��Љ�S+?�xdXпh��/׊l��|~}���	4�������OF�
�����LN��5Y/���L�q1LS^�m�i���uȺ�plDC�5A�^	�S	�SBEa����A�B���N5E"�*��D�+D�����v{�7�[]�ќOʍE7)���sF"~ڄ�*�nc.u׻�}�I���۳��M����0�0�a�_v�I9.��S����(��h�E�+�� :���Z�q���sK�� $>��'8�e&���h�r.2��|[K�9�V�'�%dև�t[�U^�K�{W�ȼ�;��rW��<Ѣq1��Hʊ�a���>��@���~�;�� ���C��8\�`�1���Q]�"i�UفZ�_�r$j��U�a��
���scu�g��mu:���|��&~�M~����9-'�
�̛�6�L8	���ϺI݂����ё2�="}����9M�H>���QX<9K"6-)))?Tq;���rN�	�?�v���Ұ�j��{��Μ@g��������p�G�:��M�"�L�F�KS>��j萇��wU���G\EC��'*��\�E�s��M�@�ghB3B4��r�]ߊ�y�Y���pl�խM�$�2�Tΐt�;�~f�qlފf�_K�ŁZ=�ܾ�8��g�����۰^e+��f���r���'_.DJ׶rز���b�˗�5c��Yx%�-n[D;�{O�CeK�[E���a�6���i����322����� �BfT$v��9��~-}�ВnؘAvנE����⁠�'5���X��ωG��x�����$̴�Ҁf�����_����ٴ�ę3--h��6�Cc�
�5�kt\��E!�a�>\��O���_�7���W"�+Ϫ�o��`��k!��#_�♥�Vb¯(^x{���K+��ڷ�s�M�*���,=k,������1�D.����v�
�'��ߍ��׏���>�&i%R!z��v)�2b$�����]��"E��b�ņ>@���}І�Wn�W��խە��
��ЍK��N���M�ز�s(C���dm{�R+XfKG�W��NK��~L�U{I�c�K�%��)���YL�Nh�B�Y	�?���V�6�sY��]�|�y�AU�^������*�1ug*���	)�.V�! kNQ|e�Лڸ��YI�[.��VJ4��T8�R�1�
��ݳ��셺��J����(�M���v��xM���.� �V�?p}P���pϲ��O����'�:�������E5��F�R�C�hׂ�ۃ��EI�9J���ݠ��(�WJ��tӂ
�m��B�7�%��P���ʫY��0��jX��q�<�
wY��ۈ�q�T�ޢ��Z� ���$>��Ԝs�dV�������!�8� ��*�I�t�Y�ۓ�N}wX�poY��+Jw�^͆é���)�8��J���>8��'ܿ���^f����!xC��n&���>��5�eç��~�F�N�Pg�]D�Xo�5�]Y,��ه�4	�%t9�j����dn޳}'xݾ��}o��l1�'s ��<h�{���]j�jN��|�Ŋ�j�[��V��=�!�'��]�#[��~����ؿ��^���I�84g2iۈ��d,��(����xȭ՟��1��"C�C�#�E>�@<�r/��ǎ1M=wD���}HȻ��/�,V��]���yOB�U�Y-60�]	}�$��d��{���/yᗕ��G��y��BgO����Qx"�sZ��;b��GO�Ġx99%�`*�N��WB/ҵ�Nn�c(�8�����Q�a˕e�4���������)����N�R� 	1�i�\�~���by(�RZ=��u�V��������(�� �=���N˦�U�&.�ױݻF���:m�s�%XIV��w���d����!Wj�0�������&5lc�o_�R�~��U^4��"��p�l�8�8�ʌYZf
�V�}�%�h�"��x�i��PE�߀$5�svW���敏�4ߍ���K�T�[�Y�&�nr=�xAj��˥r4��'��"�����$b���Q�:�_�X�fs�k��㝂c5��[ε5���N�qn�?n���G��<��;��A�`����[��4�Y�C'œ��CZ�'ZQ`5b��c�T���=���!�d)�XV��(�l��+��hQ�I�^��e�pB�#�j��.���s�~�������!.(��C�i��4n6�&D�^
$����<�+��4��^�f�� ��S˒�?�h����@�EH'�����_��ERd]v{���/̲||L���q;H���W�m��:�1B)J��:�nCGY�.obk��1��E����MB��[��-�͎k��3����e�?\�G!��q^$�������Z�w7�t�܋�i�"xr���D;@nQ���2`y s9v
� �~���,H�W)<�bl{����O�l@'��x��<�ia$�?ǢP&Gu�~��O�l���.���0�6��ʾq�\~.�����L�����f���^w�'� "�����t__<5#�PDu��:��y����ItV�~O*>��\���#y3�����P��ի��M�0S�'�G��1E��T�B��?G�=pY�Ԡ�c����\~������,`��ڙ!,���8M�%P�0������ׯ���oqQ�ԗݹ8�K�����M�{����i���q��{Eꌬ��5ekS��}{��4�^U��P�-Jƒk���FF������El�~�!TO,�$M;�=�X��׿����k�X��hsn�HA_9u���<���Ӓѭ�@�q)���o����~iuű��,N������4	!�L*�l��Y1�1�"�������kŐ�:]:�?Q\:�:x�E�_u�������}�9O^�u+�׎B�e �W�	A �� [>)�HA@g�%�I̾j��6�F�b�WJ���h�\B���'�|+f�Hk�%"��G��Ep>Ѐ�+`:���2���Q���9��ty�P᭵$3���Yx����Y�,8[q�+Gǋ�7�P
�C��Z��>�'�$w�gYV�a]��]��"~!��we1S&�Ϫ�]>,���|��dU'>x�CO���(h�^-�h�hLx�p>�^Ŋ/���hE���:���¦6f^e�Hl]�yŹ��X���a��V�fK�yFF%��pL�|�IΜ`;ٕ6�
�u�g�e#I,0ؖf�ؑ���
턳;YpO����g�`JZ\@f.
"/�u ���#�!���s2^�G��mj�b�J�*w��g[p��lI�e�]���N��h	�}2_���NLPbv���(1m���pBt�����J��X�I6�P�S���
%�?q�8�@ċ��6�A0&s�a?�wtT�?��Ҳ��4t�lP�#�]e,��t������n'?�ex�m��󇞠˓2+�3�~�F�lIZ�^UZr�b�p<(�k�������;QYJ8&�Mw��$3��@�+���x+_���,��4ߵ��n$`�Oע�xrN�%sM����|��I6�,�rb\�㫃�utt�������qH��4��٦��P�#�Q��J~�����[�C�%�=�s�^5�|?ކ�
�7L���v���	���p`��('Մ<,x͔���.�谗�r��z�Ң ���P�A<z�"Hٟ6&j�\`�3�3=4Ѽt`fVI�k�+��l�Kݕlԝ�䔓��{��6��k�3)�L�;���� YzI���®"D0&�O��2�>�Ĝ�q��[�D�eٳ��=��C\D���9�AXh���x���UϷ�8$m�L���AP��x�s���I�R$��{�h#̯B3}�j�x���|���m�{�c5��P��g�}zV=f��N���<���00ߖ�<�O�Y�-s�0�Kr:��λ��F�RU�3<��`54��O�:�:��@8��!l�[�CB�; �:IM4�2D(���	}�l�+c�#k�uE �J>�c�\K��!b[����%kyZ0���A���3(Ha�
�m�oz��M|�Oԗ��������5�7+���\@�������*�(:	ö�.�5�C���_�W����'f{�� L* Β,��^�/|2{�k����s��ɂ@G�����A���]tg?�>E�I�S
��b������>h�?t�R��쟶p/��čr]�kK���7�?$(B��nm�*�����Y����|��H��,�5��c����x\j��r�3��GwM��i��?ֳ�䫛�S!Ӑ�>>��*L��Q�h�?������o �)�F'���5��>H��*�����h�ħ��lW��QDv�y�P�3�W�֡��nN�WB�8��5S�#�����?�v��)��R��"y"��M�w^�O���Q�����{V]Q�R�y�̀��A d(E-w���(.N0�޸����N�Ɇ��m����&�``b���O��Sf�WY�0�ˆ�{Ap���Х��TH5ȁ�&��;��o�����2k�rH��������@�d.�qm=����7���G�-�D�x��ٶ���H��G�E����RD�����:�Ml�W�lCi��y�I��E �4�~i� /�`)��?�'$x�T���^�X��2�+�4�3gE�l3,��y�-.��8�p%~lb���� _4���*$���i����B�
R`8�$2*�!��Rk�仼�<{Ú7F�x�J�.��}�.#��`X�*��fc�,i0��������.��r(KI�MZnʇ ��'$X�ܾd�R �)���bW����v=KU��%J�S�gy<�����)�x8�{x9�ޚ�z,����#�Yp�FJ-���=�M���7g���C+��v,J���8~�O��]LK)t��29�"��+jV?�i�^�����<X&�齼����S�,�n�0��H����n��*�J�u�������(��4~00�R4�o[O�Ẇ"�Ⱦ���,`��Ng��s�F��$�æǼʕ����gq�Z�YǮe�:�wC���J4r�OC�O�S���q���cy[ugOIKf,ΰ�"qN\G�C���%0Xî-�0$��4#vn�yo3.qMTu�n���"/��캪����1n4���: e0�G�t����>�����4�ϧ�u+b����?%���Y5I��Ip��2��¿U��Q]�6#�_��ϐ�N�Ǝ/)IT�S���:��A��Z��P���#�
��%�����8DU�6�
�M���ud�aʀa����Y���و�D����r�N|Ou��New��U3('_ ]��(����	�;��.��ᵷ��^�,���/�6ۼ��`�
Z��c]5������pP�E�
��תϣC6�ݲrH�/V�������u�'j��m[mg��&�.ۖjݞ>?����$:�D��Zr7�����x�́w����K�M:����J��R�y��O֜6I��jF�i���/[�﬑������������p,�D�����%�֪�[��W�aÃ�G?���]-�+1����/9�
��}�}o_*��+�&2�d�oz٨h���&��s;Ra�~чI�A3�얘�N�T���v��c��E�w�z��섚��W\�"r���D��ytRyt�҅��"�\�Rj*��q�"t��������ٴ��s��u�7B�Zl��۷������Η�-���g�$����T'Hc\~���G.�Z�
�/O3��ș�
�Ip�r��ٱ 3l�ջ�/��0;������TVMi��{œ\���<==��n����fW,�[��<�_?g�r���AF\נ�rԤ��t%у�D��%I��'���*K����Q���A�	�d6�Fi3t��%����,�Xr_Qq�Tb���R�Py���c����WaG(�~���?=Z��&�1��u��;�u��'��3y{�~����%Ii�L>x
��s5��zfbi�=7���U�><��BV"�����9��ڐ�w7�~�W�����w^�/o�^Ҟ������O����8��,~�I4o8�|�#:�ƭ�eqԢ_��`N�~��p��J�͖˯J��`T��d~d?:(��e���#�P�$�Dij^S�I��6��BM��>�Pǐ�~��d�A:U%�ug�V�I�����{m;'�(�����3�K�Q��VYmH�vyׯ+�s��Fk��K�ѵװw���d��e߱�uwU�nJ�;(Q��:s]L��}�1��ՠ}�2�{�ui�������M_�I4�!=+�(6u.KpB������|F��/W�盄�8;��`Ķ�1��*���8���/�hoD���n��ޘJ��Ppi�$����~�_ME.� F��%�R�ZV���<	YU�@��bJ P�c�m�9#��^��~VA�V.�i����3Tj컜�aCB�@��r��=89�T9J�$�rM��$�}�ưf(2&����bV�|?�a��Kz@�����d�l1���&�R�y$O�y�����5ߒ��G>-[@Y��(gWgf՞^8:�7,�n6n�����+�(��_|ɔ�|ƥ�R�'�,̚����|�0h{�$)c9��M5v{f[�
���R����GTa�(���g��\C�Bv��cy���x=�I]!l��J.rte!��c��]����
w���qIv�q���P���(��W�7>v"�	��A{�WO`��Hp�۴)���"De��g�F�2G����0��m�7<�c����磑���:�^��r\*�ۇg\��q����0�sƑ7�qA�q8�������׷D*;���qXy\��/x�3m�q�"�}���8v�+��)���=�X�:Q��ͷu*Q��u۹�k\�B��pO�ShӨ��.��yꔱ� �|i���`X���x��"�?s��<�̄'���9����E#�O_��ÑM��~��2�/dk)�l�t�%P��'�1�J<ge|'��P#!j+x�'��[�i��kbs��vN�gN_�CA,����������fc�y/�c:�>��5�,U5'*�(��mk{Ii+�&`ŦfZ�G��M.�􌄕h��Z%j�?��c��R�%�gg��Ųc�@�"�J��'��F&=���nI�c}�4�b>�K�KP0�El�aS+�y��DxZ�5��u3~���
�<X��mi �z�~����ԃ����̘Ӿ ���F(1Qr���;��	�ryTJ�u��c8��i�^Gk�!�s����7|_:j�]��Њ ZK{�������<�gxD\�D�]ei/�:�)����\z��}O�ZG[���ڊ�qx$�ۛM��G���d�$k⁝1� <��D�q��/���GY���{K��UB
]�j(�����XÞ�Z�ӵ�p�B,�5p{���WJ[8Fe�Xo�8N"���~/y8���^�������?�	��og�D��c0U�a�s�O�4B��q��t��@��j��,����OW���������6M������_x�56���Ty�\`�,���_�%_sB�~�����n��xb���D�+�ݿ	N�m�[V�ya?�n�)��1����ظ�������!��crŰ�:��-�w�3A�ۨ�ǳ��Ӡ:��l�:����p-Clˌd�w>�^�7.�
b�A�H��Cg�<�U_�����֪e�"f��:����y��OC���j;4�3K���-b�T![u�0�IO����Q�����Xt�t���I�];+@�|�M�5OÔ�������)2���	��t�\$OA<Қ��s�Ǔe=IoKd��"� �h�6Dy;)nZ����@���j`�M���C��q����<x7���#�'r�7�����-��_L������f�I+Lqb��N�����(�@Xd��Bz�B��W2�p�~qh����An�|��`�N	�?K�\�r�VE�&D�H�u�U�;34���W�z���K��x���|���0�T���2���<<��m.���QGT>`U��BR@�,��~������Y<���x�����;���G*��rbH?ت�A7s�F/���?�k2��Ŗ�n�=2�4�=�uA���,`}�/�Is{���uBB�6�������"�$8�$\d�WsU埈L�?|*?���������bR�f0����qYd�����A6�����?�+��6FH���+�����t8JV�\����Yd�$Y]PDPl�;re���T�f�[�`�SȎ��ܰ�x��%a��}ݱ�w}��?��^# ��*�ڀPr�<N A5dO� &{O�"�?�}+I�.���� D���Oa�Gb3*vY�����f��#���d�E��������Ã�������n�v�5�C3A�����)?&���]po��	��,?E~��+�k�A����x��iB�A|�f�ً�$*�P8q�I�MbG��BR�(�����⺠]�K���ɼ%V,���� u�ihY7A\9:�=��&k�ͤ'����-�`�5����������3�j[=	l(�C�nI�d���+�Q��D�������˹@+�[}G�i�a��	愉_/��EǗMR��q@��(r�1�tcr6g3�ұ�֝l��1��g�H�x�m���t�,�
u'�糀�`�>�g|��I�����}cmܵ���ʟ�;|�8�5t.T�j�:�t266'�ޭ������������E�>��X>��gu�P����� (y���� U���웜�"MN�R�Sͽ?St�{t�j��j�6�'h�#��t��T@!��9�(e����F�d���}>0�'�C���(�`�0�+44�8(�6"#A�۲gm\a��P�.�d�.��H2�5�yS�q�W;���e�>�B�]�P?��Qv�)���fV����>wG^Z����q��X|ٱy鿁�X����߱�o��+�m����[t�Q��%�
����/vj']-�헤47���f��;Z$�w��s4��Z��L��ۡ�����YY[[���\R��zz�8t.�'��w������V����B� cs��c�׊
��Hw�Yhh|�� D��0��m���N�����{����}wAU��|�9��J��x¤Ԃ��k���4�=<����$���W[�5��^�?��0�ص|�(]}�e�WX�ش�5���<˂�g�1%��0��ef)�%C�P$V�53h�i����q��s<ġs?���\���6oP�$Ep�q�L�h��:��f΀蜷��Q3;��P�����Z��Y�t�
�(�~����)!;^n�5n_7�G	FW�S�=�ϋ��M��)o�b��+�[L����fcW��Rdg�=����G�7+~\}ОyT�	�P�@M�K�K��@�+��q@���Ϲ�8H��~ٲ�#�g@�"⠟��[g��`y��b��iaG@�N3mQ�,�=���N��wZ��+���O��1lh���7�Bp��߭�aCC=>P�����q����Re
�"���A<:dXߖ�zwy���A?�Z�dpȏ?϶�̴,��0��ɢlb��x���+�Q�*���>_DB�yj~cZ��N}A�Ǜ�.��;B"k^�&�(��@���d�N�b���@a1�Z���[T���I�C�8N�_��$һ�z�3/�R��)5�d���uL{��;f�Ǖ-�BL�AO��@,�&	#��������a��J>øE���pW`��h� �j�V^��e��ï�zr�WT�J�-#��g���;�"���o�xZ�O�?�>��N\��[�)�v����`L'�k�]�+��Ղ�O��-1�L�mC\�"N���"��@e���N�����t���ґ����ja�!��@��@H��.Hҝ��Tx| �K��9��G��=FJ:tXWֻ�b�pz���l��KT�%[ifz�=�X�+v�7lOv��b�kQ��

��N����x�K"�k�bo�/�
���P������ ��i�p�j�Cs\��)�4�,���xF�ODP�Ɠܭ�g{�7A�`N2��7���Vi�d)w��n��r�K��E�M�Dse�ѷH�[\�(��tXez�s�L�y)� xo����c@k��w�Տ�<#��o���=�q*�z�a��Tэ����<�H��е�` ���t�Ǜ59у�����a^F�ʟd�����x ��Y��N:r������&��s�E���U_i-��FȔ��J���bzs+4׶���1�R.}]����ǙV@��uٿ>���ɳ�ZlʯvcB��+C�6ѠWG)�(�u愰�ż��"6����W.�Tv4'#�-�Ŧ���8o	�A��
�n��Q{����A8����M��]�Z��Y�W���$�v�vk]��6Uon��`�S��PW�ϸ�s
pp��KW�����n�Ҏ�n�etww7"��Ώ#��8`�����t7��������9�y����g���Ȏ|]�V���"Z�b]��g
�����/`��PetʉsC��� ٵ,�	�$�9hogK8��-_�`���߼�8�}�N��d�z���6�ԮYΫ�KE8���̏}$��������s�J�����H�߿��G�h����#.�i���jlh�]Į����+ƌ��m7���G�ٙ������h)C�jDF\��Ԑc�����@U� -�LVv}4U/7�zORZV��H�k�7S�����P�k�M6fXb]#�d�Z�5��r��
��C���x*��
�x��,o�4vo�N,�]� ���%J�?%��7�=^ZY�?�t��H�3������ӟ	���~a���i>���{f�K�m�0L�\ �=�3w�8��;H�  ��Y`S���)�8��!W�+�#؂�cp����$E����AJr��b�>���:&���X/9 S:0�E�8p&�>;F1�`9�N��o�Χu`c���CH�P����P�%�$c���ѩ�Td}H�	�J�����V��w�x˼�

��׊�wP�eJ�[�X���ߙ�kւ���s&�T4mN��}r�P��Q���1HII)Mlh�`�o�j��q�h�)���Gy8��^���X��m�9��m?��&u�8�����t����Y&?9I�q�
�N��J���!"�����V;
�`}2y����`�S��K^+��4��=�{��������������l�6�{�2����(���b�M?y�]H���c��f���%"��p"�U:+�	�L�-�jk�)܃�0Tx�t�V�;vc�./�N�Jg�g:�oj�⍟�~H1d�KI�v��o�'�Q�6���¹����Z�[��݀'�#�2�A_Oie��@�VI3�>�*�
�����.y�́W��D�����	O�[X(�N�鞎N�P���דR�U�u�S�!�C��{�����'+����䨅�=ǫ�E��)�&�ޡ�a�҈GD����:F�]Êu*v�{n��L%���2�,%,����J��af~~��`v�A��ώ��"�u�KH(�go*�0�n���U������e׆���A��L�ߣ�*��N����g����'�N$��m$�w~���ԋ\���ɗ�_=z�J��b��W]�D��Ԃ��+U0	�'N�i�!�!nA��[1u8��Wy����,���!���й;1��Qn�>�'o��Lvi���H�f���߼�wa�ov�����u�4?W��.Iվ<EEF�?��^�5i�ۡ�y��d���QP�ɻI5�'�Z?4y(�iH};��4�e�Ju|�)��f0n�:=Ձ�pDh,�sg��L�^�ow#S__�D}����_�n�Ć�ǉ���'ɝ^MB�$'7�V���$���/	9���5�˷Cp���8J�����igș �]�� V�#c֢�:]��L��cF�����~�D��p�)>�fa)��,}�K$c&o��*�Ǐ�QQ�h�BCoG�<������sc���*�5�[�E���s�Ia!:U^����*�ޮ2��̑�V#z[_#�H6P
���$�8�1Q���e�_rԶ����Ur@p��0QZ��s��O��)�W^q���w���@�8�vNN�9�
gmE2��x�~��\u���y>'�
s��+�L�mv�@j3��~,�P�o�9a~bJϝTd1�R���<��S4i����d�e3=���w�'"����Yp���>�����c���Sb�eZu���YK�4�\8���>x�
g�=��m�'N������>�I���J�t{�K�B���>�P�cAP�/��;��o�P�rɗ�|�u��T/��tG�(��C؈�a���3�F�J�t�e��`H�v�=���e��3�L¤H�?\:�NȾ�����.Gf�>�o2T�k<;�/�1l �����Yd)���">@)`�Z��VJҌ�� ���vH��?ڸ�b���5>�u3zTW+VH��ǽ�ќ��E�@���&��ߜ7p	jcr���~s������2tK�:U80���FF���KȂ�5�	��F���B&*�i��մ�<�&����e*`��0<9��LT:}�H�f��.�HȆg$���3�^Ѫ��?���Y���m��3��l��=�~���ibV�;�����������XF����B/��	�)#���Z����Z�B�ڢ��.��ﮢ#,K�G#���$�m�zO��G"�GVQq�0ʋ�����Ce��u����],��JψO�^�L����ƀ��5(�Yˊ<���Ջz�7D[ͭ����*�j4m:��,�<22s�:�;�+&U��S��tdP�_T�o�ׁ�~?#Lb�/�:N\`3���d�	�X�!fHS�GH�޳k"��.����!���aҺ��Q����w��~�������ӊu����:�b>2"e�O�F�6C���*��|�_�6$i,f�I�ٙX�`��7]}I5Gd�l� e�-om�F|U�&�8����2@��Qޤ�%�WK�p��`|}����w�F�yŸz�����~��s�����6'�o��.��q_��<6�`r��P��aTp��c�6�x)R/)�DF�Q�mE(�☈BV�(�k��O��D���H�Yx|�_WH<��{��֤�@�g��3���r�>ql�$T�K�~����
�.v4��w)��3|�_�S���u�T�Z%���Ma�P��vyqz7by�	���HE�f�K¥� ������,�ӵ�f��l�<I��4��co��
Aed���Lx�iRK��-�nL���0_�'�o��� �z�H;��j5���:��m��·mkv�ѦT����)��TE$��6_,�;@����~h��ⱱ�fu��3i"rp���s�%�J�ߠ~��Ij�y����l���!X��+#�T=�,TX��H��͋�{����H�)!�6���?����䳨�[��s���ܤq��74��tCP��S?G)�>5D�9�)��o���׼��\���C�*��*&�?�7r�g���ޚ���������}�����I��}�6�P�@���Æ��gi��JF002?.���$��P���=>E%�8�uv�3Pa�!��{��c���Q�桤�N�=�{ ��~���[��$U<eMBa�8e�$�_
b��E��M9�"��n�l>ۯm=�]�TȨDG��"�Y��e��=�1�^A=������ٱq�읲���(3��P�۵Y��y�NL��ȱ��7�Рv@Y%��,��0�eAW����"H7{�G:�&f0z�.�6w#X�xѩ�7��2��\�CU�V��A����5�,�h<��=�p��7<�좼qE�N�3��uQ Y�D�UTԭ��8��
)��8�5�������9�iS�F�wQMr���ǿ ���r�$π���λ���#@��g02j�[z�D�&FY���쩇����0g�"���ޏ4)�l����*"XiIP� �PB"45���^GӾ`A�|���a�x�dT�<��GT��*��J��DT��wI�K
����$��Q[$�7��	�kA��I���T��NTz	��m{)����~�Qf�?g����Ҵ�\��#7�Z_0Pҥy�=��eҀ����*��.E�X�.s��Z�A�xC7]��~��J*�Ie������!{����S�ak2n���j��%�^B��$+ߺ����,x�k'��Ѧ�?�@T��F�x�fD�Ƀg~g�}�՞�ѱ����)C��X�ܧ{�4���?ő�,9b&R�'};��n�W�#��?
�Ӗ{�nN�o�n�9����.#�+�8S�ه(�;�]����] �;�A��JEť�W�7d9��� �^ˍ����_9BM�I�f�|�*m�6�Q��S2�_�p��$gpі{�ڻ�C"q?�l~�W�B�����fWO�_Ҹ�D!_�g3%���}'�?���s�U��8#ʙ�D�VPP'��L~(�$	sl��W��! ������y�W��� g�����!u	���L;o�b|%�+R��5�:p�c�9^���e������C���Rpĳ��2���G��I��Ȼ�?�Qw��M�˥Q�y�r�a�)��5.>kV<�:q,S'�S"��d�����v��։e{�cB�g:i�|dטڵ���ጨ{�x<g��_�i����);N^�d9�$U�E[B���I��P|���h".'���՟d�o��ŖF�Ļғ
�HBԛ�|:���C�w�%����a�n����*��V��v��P[Z^��\٘o4�ף^��\8�Uz����UE�7{�� ���{�PNL"ޡ����
�(�VS��
�L�����{,�$�D%�d�5g�Ŭ�V������j�<E�wuk��Bbx�V��P��1�>�)�[�Y7K��x�Ls">�� �&�d˟r���b<�ޣ=��cv�M�X\�2��q�i��)��[~�7��hU�I�Q������*R��@�r� v�9��\@����Wk2�UG�ɷZy��U�nHO���2��MB�@��N�]����^�ޞ��̴�ܙ��S�U���`����I�*��_I�}Էw(�M��0�Š�Q_����Z�t����wl�ǅ^V��(����y$�×��𷦻Ev��yl+,v)x(>�SWV�u�<i�x��i+̰���sM�necco�w$�����Kۤd���x�
���ME�u����.����e�X`��� ���>M��<�N좖6��/����퉤�DtP1p��6�L����IpOm�� y�Z��F-�B�Ď��bb�o
K���0�����ơV"6�XR��q����P��
Neϸ�Y��I�>P��	��\l��q���󛓪���A��G��?���mN�#B�+��+�SQ�'�AQ�m�rX��q<�1�����ks\�ٳ2�-��#{X��@B��-�������W4������ۯ�$�v ҿ���ddW�I$�[�')V�D�	o�/тD�@��g�q��F:qɏ[uH���}����C�\{�oLк���H�-R����$��RSi�u�� y\�ɯ��mAzs�bȝ�d��ޕ�z�R�ӞSԿ�~�+�E�|<�z�s)������>��qM�;99�t��mQ��J^-������v��͌��T�3� �x]�L9�a&R��|�������m-��,n���J���_�7��*J���K���[
���(۫��)b�+��oS%frR+���=Ld�o"�~�)\�'�|����M!�ѳ�m[�z��:q�@�3�NHU��ó��t���j��=Z7���R��U���X��yF$����8�A�o��� �T!�w�nv�<��tzM���Ȅ%��U`!�O�7����������۾�=��M�����iq@�g7��H�B9H��$-����p#�q�?L	�^+}�	ۘ�=�*ED��5TN��p+���$B ���"�O�����Q�Jl�$����O�J]U#� ��1=88X^���N���[�8�b���Q��֥�g��P�χ^�x���������9e�
T���5L��9�wӢU�oi'	6C�	���g������/���6N +�./ٿ��P'6?���3�����ġ�TP�ko�j6��� :��ۭ�d�Qww�O.�s;�*���h��d�B��=���fk�Ƌ2o�'��}Vˢ�ߣ
rz��Nf+�h:��>�\9QN�ݦO���Y،M�_ˬјdν7�B�(L4,��o�aOO4Q�NO���G�$QwAO�D
��7��������+~���M��
5��F�}�f�*.zG#�#2�����[:ί�߿��<�DB/)����QMY@į�jU1�|T�֢���0}�6�ZM���_�)+3��@,�ʛ��ig_b)$�ǋ�����¢��ے�I����F�
I�<J]����[!ԴkU�tkw~���$�����o2�v���>�����5d�o�m��k� 9��< >A)&&�0���.z��*�+[�8��<�{5I\� [d���`K��&�m�,��让�����ӳ�@��L����U��4�d�f�}�,;�ڌ�\;�������>z��RZ��*��E��I�D�5((H�(Z&�8�E6�qU\�w�|�m4����W�2Tg�af�y��7N�/� +kwA�AO�+�\��M���(~�\�p�xq?����8��y��p9�����[����3أR�q���M��Ӿ_�M��o
J2wz5ʹ?G��iQbOO/2VK��=Y�tc�=<�z4"@�\�키���{��=����6��H�HQ�2l�2 u��5�ʉs��.����M��DEr8�B�'$$&��kOdҰM� QVJ���#��6��-�X��i���	A	�(��d��.oyC��Cs�>�@$�='��m&�9$����X�l������TR[נ�N��s���-�sNG��� ����\h˔���w���f�,fڀ�O�u��$��!�eo6�=��6�ᠹVW����ƍ�M��
N�l�}�wK�i,L!:\U*<W�|��~��kz݉f�h�M�o�K����9�R:pX������j��_۲P�o���}M5�I����򳽪W8�X�8�-��MT� �Ȯ���9+�z�WA������]��L�J�͐;%�����:0YgN�&!%7��!�>F?Z���W���KeV��;�)Ǹ<�&�m������B��@���TV`��������[�������ʘfU�$��򺙭3w �YݧF���SN��v����.��>��h9t�P�
�ca��=�[�N���G�	ѩ���_M�_������d�o��\�������76�+��V-����E���?�#��3Y@]*P��[ؚJ0�-�K����/��Y.wqU��ױ?��NXRw�~M	���I�Θ�JNr���Ͽ����c0\�so�3�9y��[���/rr�������w�xqj���C�O����,w��i����6�H���_{rȱw����� �nc>��88���P���Z�i�amM�@-�y@���m�d�	2ۻ0a�llC]�\��۰���u�w�WQOW�{UU�u|��z)[\�@�*?X&��	��W}�v&M�}0�Z�wuEj�� #���$�҈���M�n}k2o��3_[�k�b�o��u�����^��A^6��d�W�Nm4�jT�F�3�Cz�}kZ��-�<]�O��G�n����ۘ�/6�ξnf�8��k[Ī�I��<��L #㴓|�P�^��O�W���I"`&h���-��z�%���G�Ðb���m	�)�e�4Y��3�ub�vX���?�y��+^�M`P���ZUxM�g����5qH��RDe,��A��'��Dޚ����n��wŹ�s��u&]$7C���]����P�H	��{�S��w���=D����y.�ŋ8r��_)#�<EzEr���w�!A�S��M�9˕{��E�l��Z�N�G�k!�!�4��o�{�y'��1��݄��A��b�&tO�%E�%�b�9%1E�������)a��?Z��e~�	�=X�Sj�X��$I�ڭ7�>�l�@z�ᖕ�����ti,s	��/���M��
ż���X���"^�Z����$
�h*�z� �PB\���)Bq��/��o'8Q�|��H>t5�$#~�t�X��Q	���(�����D\B;C!����>J0�300�8-�Xu�����e��^�/���Ý�߳�S���R�>����U��oV#J��N��ڤ@��I�H��i�P�!�;��YĽ
���k�^Ԇ��)��ޅ���O�E��a?W��o�=0��b(�-x��őA�7�5S����v�[0蠃��G	������#�l hx�Z���E���m���-2Ѫ[��ӞMP� �ږ�,�Cζ�N���K;�!���CYy�H7c]�L����1�"�������=��52���f����M��t}e#L�O�P39 �'����:�\+��҉{	XAG��c�s"��O�� �;A���Cg�t qPG7�Z��7R�|P����Z�(?��|���sMEE������	)�L�)F�F�%��`".%e�����'**c�6��W���T�?�=��F�'2�@�fM����WĭwP�Dp�jz�
L����N@�?(i�>����`o��󛵽��1����{�ːf�a�y��J����k��g"Vl�i�|�1��� ��?(S������i9n��0pԎ&��>s�Ti8��_�W�\�G�Cs���F0��ѩ9;�5���:p��d�Ic#���%dN��I�
���_���;�
����e	�	��惭ڎ/��b��g�g�@��u���0(��r������X�����mC9 �������%���g�7�����0?\Knu� Q)�q��9�Cƹjُ�m�9Zy����GL@j�	�ՠn7�[�ey"s,�H��>i�dU�;��Rݐ֋ʁ.�U�Ŷ��� �	�QϦD!+iF�z��qN�,����\�H�K&]êxsK�3��f���)5����:�7f�~Vѯ͉#}[�-�Z�ͨ�+���'BTjx�P����� �����!�b&�2�N�1�T��'�����'�Q��;��\VÃL��ldڔ$Ǉ"���m��t�4���<x�'Q V�z��������A�i�{�ǀ|�5h�T �]��	��V��%ۂĘ6d��<��i�L�')��R
b�wt��d��k��=�/2ȥav��h�w����쳼*��q�(J�+��R��A�I$�-�-���DI�;��o�qW�k,*=h'<��(k�;[	<����T'�	��P���&�Du�V�vs��?��J�� ĎpTՏo_��u��?X=��O�y�,g�C7�y	�@J����e��؊�	ךZG�Sx�T��"=y�� �L�`�>[�鰳�_aյ���������Q����իA I��Ť����m~�?�i�a�NN̪5/�x�ۃ�_D�:�ؑvu�P2"��\��VHrqn��,�ώ	��I������7Ǝe������M"����Bq�d�ܹ l�rf"�K!U�99Ͼ;���S�X�C�l �WW�V傁�|��g�zOى���ԯ�6���+
x� �@ �Y�3�c�	���9���"8����͇l�ilU�S������ �������
�)пݻ�_
IrK��bΕj��o��/Z��Z���I��o�F�����|7�'�UyA���>O��l<�	ZQӶ*3->5��iRw2hV��M[�,^���ͧ _�T�w|=G������>q�����RÆ�K��@� ��6e��v����qv$�s�1���re�U؏��W�����i����~~*1�>/���v";��V�t��EJw|%Mƽˮ��yu���N��7�8�M��,�-���������$�������}ca\����}+J"������TY�� ���u��uO w�F*D����:00��HR9c� ��)�L��/.�,��* �D�J��������u�����o�Q�͐}]�67G�
�y}��~^
H��,�wmV@A��e���t�g�{�R5��i	�v�������l1.�*�؍ȆQ�8kh�W|�1���ε��]9#�*g��}�
/���t�qGw<T`:l�/���3���T�4.� ��>��³��UY�i	�8�ڏpр�}z#_��_3�s��=+S��h�;D���~tt�l������wD(����/� "U����a���'�挆�c�.�Fp��~�:�	�L�{ۮ����� NOb-� ���%��ɸ:�+���[9ڍ>���(XN>�;�ҹ{����d�'�S�p$*�>7�=�g�Z(^
p������KT?���8XEAf\f���XU�o�R/�
42*zc�kCF�����3EW�m���yD[z�n"%�AT�����Z���/�r�/M_��]��C�ww\s]:�z����a�uu�{<ܖ���WC�c �l�
����5�����'xp����|E���ш`t:H�'���j���7�x6�e�RC��w�nO4Z���4�����@�`��ց��.u��T*���(�=,��������|1/��A��,r����ˊ�A��y6xD�̡����=���7�B��m��u6���@�}ۍ�Ǽ�_�������>�>K���_	vR\ FW ΛK6r#w;!�g5޸:=�����܇�5�s؉�6C�Zִ�=_18j�B ���X}j��� L^�:Z,8��ި4��?.�dδ����)Vw�Ī���g�U`bD��Cl��	#u�l��=�
�^�5ѣ��>�7 &0Ѝ���qi�s�?4�=�v���ˢ��b����a�tm~�:_{'VN��r=�lV���� V'��t�0����yW\>�ڸ��<^ӌ:���D<x몤��"�^ẕg�)���A�`��z��������!:N�u2�����l�����ܟX�{b�+�
�	>j�o����&U�+'�T�m��0᥄)@���t�	lZY�؉��y���3��o�t�\�fԴ�+Jc�����:�JC�C�4�d��0�W��>�q�I1�o�m��6��Yd�d�ns���R��&��6#��σ�uEV+ {;�mZ���� �;�JI�񐞝��oĤ�h��=�E��-�a]'�2׈5E[��EvL}�d��6�������?��-�\��ӝ�����9g��^���\&{J����WXBO1@D7���n2���h3DU�U����'D��ML��#<e��~'�{���U�Y����������!;��3̄�Q��^|G����	��0;+8���OD�+���� �����������S'�K�V�k���?&�d�;�T)?�?<	�xj�h�=kb[�
�ZxS�`%��4G_�H�O��,.~�eD��^��a�,'Lw�2�講�g���q���7t=����܁���7�Y'�����H��{���n$[\a�
�J�kf�b��g:9�C�$��Iܗ�a��Sy��K.j����u-_�-F���r��Z�ا��cz��JV���g���u\�w"F���8�Lu�ˇ��6��������;���I�#�S{,Aq�}djqu��h��F��V�[
�[�*?��FR�ݫM�s�z�ª�xax�dH�����>V{#��<�<^_�Cr�����1ӂ���{;����ɣ�������5�5�3k�����6H����ז�+N�+6�8�F�!P�C��Ҳ�o�񞊺�&P�<T&�!S����,���֭¤z������ǧ|�[�?�X��)*�+b�-��@h8,�ŭ��8Mt����C��P�}�[��yDCtw��r���|���%aқ�$�BC��^�	b˴�,�y��4kD0B�u�o=Ɣ�T�$��0E��sHGޛ�O��p�뫆"�tC4f��dFN��]����F6Vv��q����l����l���i-�h�������BVy���af�,���*+Y���[�yж��1�3�&�~im�w �����(����KU�̟� �2���l��>RR��m��������֯�id:9%�\^�]�TB3�P��}�tz|O�Y��n��le�u�)�9����A\(��/N��fsꕬ^Z�?azB��*<ǃ?�}<y_�[ZJ��h�SW���}�6�$k�Ƙ��ȹ�V%79 ����G�V��
��t�1��L�89s��7��R�7;��i&�A
�����b���p۾�v}���̓�^^����=����ώ���sh%z����g��K>`L�N�o�����;�D���� c�(�9�X�8�<pSM�_	#W����&3\F���iE�wm38Xڲ$�����1�<�=%O�N�KWyXKSP�Y���E��Ļ�!�]�'l�];=���R��-�v����0��O�� ,=��-�^���I(��îG�z�<�Ӵ��2�Ὃ��ܯ��:�"�uB#����}�gw_th�����I��)�� Hp6�U��D��4��)�G�˞[�S��T�8�{��sS��an�£�Ǉa���%)��^���do�G��� �������kx��AuN'_C�����Y*�2��$�g�w��/1��@���5h+1�0���tw����OHn/]���������86R�f.0�h�,��o��$~�7W���Ww`��ɧ�Y�=���$)����r���.i#��:�����~3f	S-�D�U�:s�����Z2��;tz�����N�����m���_��P��쎌���'5a�8��{e�I��������z���+�Q�/6s�{ \ԩ�Zڹs}'p�������/0>�[�oˇ�Q�E_ǏCeܑ(h�1�U���L(7^�CpXT|bdN�'����?�"���z���ó3g�/{�K�@tk�5�I�����L��/i�j�S,�f��'Ȝ?�*$q��-ř���b\K{�-�Mj �50� � �y�|�Z�"�̌炙���t��Kr�v����&>m�qrV/�E�|��8x�K�˙��d�]ˢg��ߢ����x�q�#Y��E��!G�W�E�0��mv�����*J���G�WB^\����8K"e|Z=��E9$m�o^4�ɔ1������=��kPڽ�w����\�!o�� �
{���<x&ۿ~��V���_/��?��� r�C.k
�xjy��&y�7H%�W�$��������mј��-��$�"&_-���5���S�DD|�8v=�ʭ(=<��U�Q���w����fd<e/���E�log�<|n���pG�L_X1�?,��ҺrT�C3�am	��4�{�Y�F�<ӳ#�)x�Q@�Q`��<��t^-�,cc���������W���Lx/ #��C�ɔ�'���,0�'�����I^���ɧ��n=�yhE���$�q6��q\tC�l�w(��E��s >"%^��Ûp��u�K;ago�^�d�e�%l�$?nvv��L�<1G���n�?�;*������K�w<�5��L`r�	�~ZԱ��Ƞ-�߾'��Lĸ.
Sz������0�{~{��aK�!�T;���;��� �s��H��:�`���ʥ^|\���p�A��ǲeR\[�9ͣ-#p<a=��9�h���n�O�O�̬�}�Ut���A�]��[k���;�]�OS�����A,69N45��þ_�M�7�����7M_z����f��{��Vl�DԻ�0�s�~:�9��hFM�	�o,�T+�G�4�����V���^��Z�Vp�Ԯ]�J���^�Jס�����7�{�9�i$�xbv��#d]nI��5�z�ض�e�:��c5���|�Ѧȁ� ��+��7/���է�ЩP�k����U6I��ej�	���.�R�3��I��oS@l�gzʏ�����m����z��Hp�g�e����d�Z:��O���Dw�/����ϲ�x�EO�vT�|3X,��yk�C�$��y �A���eg>��=̱�Fa��.n2�#�����D�ߜժ��9��߷[��@�1{	5Hڳ�!z�.�$>lR�f�y�մ�Z� }G����
�L���V��A-@ΓS��Y��k�[�=FV>���i���i��Y�t�쩆��]�t~�!ci���,Э�D�9'�y٠{V��@��)��$���]{��]�v���%N������)}q�p�_����e��M#����t5��}�{΃��y�I~Mo����#��5��:�h�y�#k��m��.�)���37t�pkJ�����K��l�D�i��4�NU~]E*�~fF���݁�;�M����k��Q��Z�E�r&;=������n� �"vy�G�q8Si�b/����;$d�5 Յ��`Dϣ@�/��xd������t� 3-�R7��`�AS��:V���/ܚ��5����֗D���g���J���ws��ux�Q~����Ba`��j��e<h��}�,���ٛ�p�݇^mX�T�]cSf���~ڶ�|�(�Hm�ࠒφ�6����)�3ϦS�#��r�.��\V�Tā������~��W�$$$�E!w�D�r8��q��F�3d6Q<:��G����+�Y����b+���	��U��\Cو ��Ub���V�C"�P*[�\���V"�4m������lq�]R��/�����e=����Q�E6� +�'^����)e���b ťCE����0�2��N��P��Ӎ^�%U�Yrt�+�[�����	�o<n���W�~����MD�6�9n�4�0f����(g7z&C������{�FC�q>ߘgv���C9)|���Q L�3�Q��sS����z���p��&G�����&��I�i~�>Ԟ�Cu��@���ɳ"���?g'�
���ۯ>AVH�߷Y늋�r�:¿c~hnJ']��S7{�y\n��|�eJ�/R����ۿ��oZ���%!�C?-�@>G��,sz��]��[;Ǚ��k�Y��)�
ح2٠�i`K*���]�4x�R;��B�Ln�f|��옺��(��	����{�yJ&K|�N����Y��T'��Mj'����󮛇8�Vw��Bz�psU/��̧ՕW�e�Q��A�Hy����M	x���%f��t6[��xs�y �֫�7c�G��BdY�Mj cM!W��$�v-� __���/&ف���S�x�z<i1V�>�h���������SB`�(��o>�A`����������ζ��}ܸ��8p����zy��󏖽n6��z�BIZ�7�� ��`��5�zHE��$�4��Yr�'�Ρ�J���Ja�g�~�U�QT��=�[t��4��{����k��/$4l��:=��|���^3�|L�����@WM��� öeO��>����.���`Z$��ks�k�q��5�-8�f�Q������;$�>�o/}�S��H���r��Њ<�׿�>����)50�N?�~Vt��e�S���.�b'M��?>�^������g��Ӥ�+]BR���j�jH3_����X+�:���;M�n"���>�,1&]�>MU���{ήr���Xi���1JSB���U�����	ĊZ~�I�\���X�\!�+|�W�]���KEHBJ��v�vxf9[����� c��!���L6��m�U���b�NS�X+�Ҁ���Á<��Y|�r��<�B�%�;D2�:e{L�o�]gIg!z{��p���Ҹ���џRE��%T�q۸Dtc�x�D.��N)�e
�"k�S�lS��O����, {��0���&u;�A��Q�k���$u��mF=�ȧ���OX��D�T}+Ԍ�̲���A ��8���P(�;*��ݍ8Y��8 �fQՊ����6��w�W�10��M�~��Q��ߕ�(v�!++Z�j�y�buk28�-^%h^�T�����󠑤�N��e���e_�������U:x�M���z�����3L��T��Tǻ������oy���=�V�A�zc���A7�9��I%�Re X�и�K������yx˟��Q:�y]�(�y�`vq����� uT�%]�ʱk����_Gbc�V������B�an�Y��Ơ6�� GsŚgQ�c���չ�
kȽ���͗zì�UނS�p��\M�1^h��k�;^�l��>���0�+-QE��ٴ���T�{���|�>�=A�3=� �$I���9І�m��vR��&1A�zrkf��0ЌϴL|%H=��d����`���ο\g�3����O�W�ݺ����i�+�(���v-,���M��oM5�A�ə�!�d���:
��/S��zza9�N�&E�2���?����dgv,��K�p��@yyy�Գ�E�V޾�C�����O��S"�0:�4�@SW�9�S�&HK�˞��4X��G�_�)�*��IIsá����{��><ߛR�n���y����|K��]Q���Q��]_��C���>a#ZH1J����+�쇭�XT�8h���H���EO8+�>'-T�9��X��d&��'8S�W�yg@�]����]��qyMi0��o�W��9~��-�����Ϙ��A4�yހ*,�v{�1�i�Ub��گd�7ʪ�����}��T�H�H;�z�����9F�c������,�"�۳�Cږ��A���SNT����(��K�֋@=�q������B�_5�-�J-��?�ќTkhV�R��*�hc����$.ĚL>�tz��:Z��{�)l`Ѥ�.Y���E)5�r�D���e@�]�_D	AJJ��=@���nP���� 5`��@R:&Fww�;���>���9��v��㑧�L�i�O����+b���hn͢�{Eai�Gm�(;Xm졶_ ���F7~�'ݱ�=Wg�bUVWΔ��������a�k�J�b	RP�0?à%٘eЗ\�ɳ��\��.���
՛�6�N=(~>3y�.�ʈ=YD]�ؤ����9I���e�;��v-�+��v�V�3k�w��~(ש^��^^�P�mԍ�Ye�/��������Ķ�����2��Y=��j��"Z,��?��Y|�}��b��*���A���A���׈�߾�U�sSJ��tpe�'#c�$3b�H*�l����8�M��ʮ�ʲ="�D�.������,]�S�������FiO�,��{p���ŧ��=�R*[yt!�f5�[��*L��S��,��U--��#v)nҗ�2��
�D�Ou����tЊ�
�4�y_�ٱ:�j +����;�����%ׯ_?���zݾ���t[�_3M4m��?G��X���nD y�^n�9�[{�5�@�����$��
5����\�3��N�#<v����ս�Ox��_��[9Ӫǥ�0j�?8`�3��E��1n}^�}�(����:��8�*TUk@ k�*b�x�nB�ӓ��]7�\���j�x$�i*���Z�4�U`���:'�����*����K`�)��!íU<�zE�h����[�~C����I^ڐ2ǫ�ם��hz+�O��Ou��� ���EgJ�qq�R^�E� �=KSϩ��3�j�s%[�J�z�a'��4X�tt�CN�7��Vyf�8~N)Q��z����cW b� ���_T{Ӿ0����+���ñ�ؓP�,mAYy�^��������� 8[페o���t���l�{��gR�CE��Ag{p�W;_t��1f�r�c�5�ʏq&1Gݲ���ق��0���l�y�S��h�i���NEz���%�1&��3Yq� w�i���S�&�?��U#�;GYv2���ı��ѓpA�h�ǓOC��!)Jl�R�
�9������+���N�NO5�4��E�;��	��^AE�R�3�E�vK�}%8�B�����Ć�ow��v81$p�-M����kU#�{]�\������> �X��%˰%�M�@5�
�*ʒ�{4� L��֫�M"8϶͵ E+)):^<��	N��ėn�F,����*�3h��-��U��B"!�M�����Y���ǳ8Vj��gx\\����Lp'���Ţ����r��s����z�mл�T�������c�O}���_S"�5��]B*���]�)�@�h��FEi>�$lM���#x�>f�����*�O��z8$nbvw�#U_�5�?���R�JWL�h�kȺgܥ{|��n���1O����9-�z���w�.��UvՍ�,�����3﫪��
U��'t)wz?2B�9�a�>��{�V����9�9���m�Q��
�	��-�I�e�	2=.]>-��>�]�fx�~Ws6~�2��UUU^;4?[�? =L[n��`�]�Q$�h'.��s��^���C�)�[�/�&��b'�B��3�j��25�pޡ�˲���?����O/*��+�D��Z��|y\��_>9oa��;:a�bb�����q%�OHH�Yڻ�%����'v����{�kmOB��_��
שv}Z�49�)o6�|�_㵉�
Kĵ�X�<��rR��z��+H�!�{1n��1�RAo/FU"1��r@	�L�9����f�n#���󃠨�LH ��z��vcR�>}�k �,��Ґ3�ԝߵ�^x<"Ӽ�9�]��:;/�қ��������U5O�##-z�C�$���!��b�3��_�pXƮ���ԆO�N��ɀL'�t?SYۏ4:��F�򦑤ej�_MO�������0���h�U�+�5֘��
L����j�9�%0�J[`O�,��K�m&�������?{}�b0	pM/�����ߟ�O\��aGnl��xq��:��t��<���}��x�G4�i���P�U[�qZe�6�tt0J[`�d@q�<���]�\P5Ϗ1������#����'@Cqh�y?]���GQOUʄ>%��W^9�+��<UķaI��_��-Llյ�v����\ZP�4�<����S˂e6>����u��Q
֭u>#σ����>V`����A^{s��-��-�>��3�~I�R�D߈ٸ��� f	�=]��e���
��z��:kY�Lo�e��U��L^D:4A1�V).�811���M��],)N9�"o/&G��$L��~E��v�v�q8�����rfPϧx��G�&?F׮l�I�.p���� .�~*㵒��W�U2�h�S��N|��7�]��$4/WWq$Q���Ӊ>��{>�@��y�D,6Y��AS�Y8;��#0�g���B_^6��1]�Y�?��$��8?�/5vm*�f��e�퍴k�Qg�	���.ˡz(xL-�p��e߻��P�i��w��ݪ��{$��q��Kk�4:�����7��gO�/��BS�xہ��*�Vrp�I��^d�nĳ�[�w�%0�K�i���rx����ydrX��?�~�z���*��}1S��ś��A�6�cJ0K�U՚ 'G��ջ��"7#����]����3a�����]�-"Z���#!�w��p�h��]��
�i&�M �U��*��2�:_<���1�e���6B�Q���1���s�����jcn2�	g�*a"D'71�U����X�f��&�X҃�9q<+��~����Z �Ι�ܽL)�nD�z\G��������aH�c����1�y�%���N5Ûş�}}D�ƽ¬� ���w>�4ː��v�0��}9�0mA��/��
[�ْ�ӆp��ka~�[]X��it��y<	hؘ�.��
�(Ҡ�8�U<`��>E�����]~u��6��9�`���id�PW�F�ԶҲ3P�a�{��ws{'�!�ߩ�mH�ᅳ밝�51(I	h���G[%Z����/ �2�U'�{,8�����1�4��zހzV�s ���h�En����P�$�bh����R�Ȳ�s{�5±pp�����b�=`��pe�B֓���r�1�M�*�l� )k��m�0K]��$�!v��}\��W�`L����[��9Ͳ���_�:WQT�D��{|(����@�N��½�����Qp2�̔�Q/�,���VչO�yt��,��9��M�@j۾e_ I��1�+b���Y�)O&�tW5单�ǝ�7�J���"(�zғ| �Bx����|f�Dqj9o���<䵕x�� JcI�nD�͸���+��a�<��]��`� uhK|̱wz�g��O�WW׿랔o�PD� �yp>�e��E̳��)`�܎�'t1!Q�'61`��e*�����A�h{Z�)j��~b跤"�V��!��I3dZ���jJV��OF��Z��\D�:]lU�Ϲ���]`��Y��|���Ɔ�=e���̮�)������ש+�%�ޢT�'�I�s�C��Zlll�:��θ���us+]�G��`;H[.�B`P�a��`z�yg�*�]����d�(��`�H�������}���\;}�Tr*����-2XJޜ�=������Z����|n��?8���s�!�����7G�s��j��W��H ;�v� [jU�`^�]����6�_��ۤ�V�J@����ፅ y��Q�Y^���Y�<"��#�<�pq�"ިb�|���VQm��ǥ4�c�7R4� (�R�2�+~���Բ�c�F�E���S>|�4���p�������O�:����qDe��fPL�0(��i�ewyci��r��K����~������Ns�����짚I��+�rD��e��M:4�N/��I>"�	���bx�1��s�m<�"*�"��n�&�y���IBo�f�9��HK>��4�aei����x8C���S��M=<�=n+��i�W��hl�۟�q6�^e�3���h�[����i��ܸ��Ώ�+{�[;;??o���H�2S2m_��f�aB�K����'k82Y�p�j�d�9�[�(���bW��u�@�������\W���\��r1�����|!G���Ӻ���}��xh4*������p�^�v�	j�1���Ha�v�;o���� *����'Ӡ�ۂw�]Ԗu�'{�/�,���J\o�a����Bk[[��l�:$b�m��`�ܽ�x�gG}ڝK�?��֘�u-����|�L��rZXY`/���_~��%�Xbn�`-xjH�x
�.\��8�>O36�C���v.2�E9-;V�euLm����G�{�����&�$�j������4�����"����Ha?R�cO�(����XWC�����TK�jM��s�1��!��E�-�8?�\��U=�s8�i�1����Z�i
W#�N����WWiDe�Z�|�L![��uw���֐��c����b����浫+⠶���Q�p��ͽ��qہ�S��\�����4������n*�cBP]������Z��G�������PN���#�'R:���-/;�@��<T��h���U<Յ��z����BG`޸m�p�)���]殛���q10�#0�ţ���6�0[u�p��IJpU���S���Ŗ�n\�۳W��i�%�l��z�ٻR����܄kJ@����G����l4T�B����M��[٧��ą��SsnCnB��ΰ���_�������fb=��/�ᾣ�/���jjZ��i�$�'��^s���S`�"w�$�9���d3Y�/_^�P��
5�	}2�38^��D�dY7�����pu���!?Iu���Y�j�W��x�[�w�J���7�����RT�m =���y=?�n��"��09��]�Ll9���:�SLD�2�x�EmS ;��^黝^��J2�Ӆ��z�]����������+탬|�Z�IB�,'�Rn��ϓSm�eB���Ajg!��0/�u��@�0�^5�iGr��$���1������������>]��7�x��5�cVY\��/�9S����]���%�2US����T���ߕ����,��[�M��i������Ǩp~��a����Q_���&�t�������ٙB����'��$���:BEހ#ؗBGnlC��t4���w�_��D�mڻǃu�Z(� ���=����:*4O�=���~��u�`r����o�~qn3���EF��R���Z��6�?g�C���}���>Ԗ���N����y[��P�9��֯>��Jgm��}Ҋr��#�B�ዱ�b�GG��&,�b�lƕ�˨����F���k�PI*�~�q�sa�T�/"w{w�@^g\��N�w���m��"����H����f!u+b]7�z}d4Tk
�(U�O��[���L�E7?3-bM�^��^�ǜ��Z�H8�q��d��/X	��!"���.�k��'za����y��v��r]
IB ��}@R�0m�֯ Sm��P�9�ť[�1�ͳ5uI!�Ϥ����)�Lr�����*����ǻ4�������f�C�8�l\���{8�݆֕Luįs��B�?�ˋ.3G�5�?w��@���0����6�y������r�~�A�o��T�L�'.���:,��^ Z9�9|�/�-��
�PK����ģ%X����u	�D�jI=5���s�	�\I_�O�����MW�`�dL�b�����e�C����{��bN;�H���s�Z��k`¸m�fs�6'uqa�;��dȰOq�������n�J��;�����'��C]v�Ɨ��^<��ڂ�г�N����3�V��[�Ʒ�mkW[ d����/Fh�ϣwm(�b�Ih�<��Ġ���uuj�<ť#�9*�������9P����B�Q��C�@�FG��4>?��G�x3�F5�d$4f<j&��+��]\����ެc�/;lk�D�=�nnM��ڸ��7��Z@c��{%}`G��������'σ룴�t�*}��s ���-V&����@�J�y2Su���^ǩ+m7c(��6ҊCٍ�?�?<�>t>���v���t�\�R�U�?��S���r��$F�)i$���OBb&k7h�6J�N5Jo���5�}�?�cO�L辗�pe�岪CA�2�v]� A$휉V>��o:kӘ�j�p��T_G�n�D���Q^�6�}v~*<)|D%sE�:�����Ml:�]���g�a�}`2�D����~<�g(Z���&��T3���g�)/w.,� ����]]�!վ1�c�X����Ы��=$�{�Q1)��U֚fw&��F)�4j�֬�G��I��_�1'4��N�O�~g������T �9��<����o���􂿼Z�
U_�N_�&[`V��>ǿ���%I>�.��j�+F���O��,阄�.������e���s�L.
���47�
�J����H�������� 7E��MaK��,�K�a@����Db����fH�//_t�!�
ˏ��F6�1@��Z��u�2~��^&�c��I�|մ�K��F��ޣ���?ưXc
��Y�i"d"*��`�߆����7��A�v���+/'yHK]\c��%�F�?�}i0׻��mܮ5��ej�qp+a�����o�~+�]_��qB�_�e'�<�'��o����(�]�r���W��m��l|��|�&K��G����r��Dl3$���do�md��CkEV��f��ޒ�2-܇����>���	���Sm�p=+^y�&��8M���h�}�aq��(W�?�jY�db��@�DP��w�ǉ$'�1�/�܇}�=�7��B�	]\�hw�^����t���I��z���ʵ�)���hz	��{@a��i::m�	�1
3�R���d�)�Z��Y��ۣ�1ҮC�[��?�K�ɡ8�>8�E'vӅ\3w��*3�࢜�\��x����j��r�hC��Jڤ�Gmt [{IR��+�wR��	�Ow����&���
��A�g��@���w�e��4#�0�ܙc�Z�x=�{��,킨sf�Ū��K�4(���srg�R��nZ�'�tG����\)?� DŎ=R�FɌ,P���]��=K��'��W���9Y�׹��Е/��iY�V�#�.X9z�����Sպʄ:�^!��bG��b��ǜ�����F#�Vc���Iy��׻�NY�|��wf�v�$���|�����ɓ���/j�DLo6��l��<��2�k߮�*�n8�W��:ZX]E��\��&�&	�+��4���$�5K$�Pa�x\�(X��4e^��,_�b|h(*�B�	��i��P����0�翉-�2�+�`����x�I\��>�ޙ6��x���!�j�����a�w��2莍��?�
�}���JH�c��Hm6�7G������Ԫ��I��R���_=<�3�� �W�-��aШB�oe�\)�㜴*�& �F�կLy�(.�mbo��� ��|�C��V�e_��H�u!1�����\�)M���̖?�u�=E(T�B���8��
�&��C�-��t� ���� vbd򇛍׻C����X�@�g;��+:�w�
�߮���F^�,��+��X4.ەo8�l��{M���rzg��5����Ű�m���J(WQ��u|5e��-'��C�YN��剜|���ϫb�&&�9�~YR4���~~��h�@7��B�9Zc7G��G�"����W��郖C~A�s�4z����l�ѴH�ns YB�B+�z�ya��4��Խ���H�!��^������ۥ��CG��L�_���	;�{p���եM��'�&�J��Lha�Ē�����$�W�'rx>�Y��/!^�n�Z�+ut�r���=�c6^��9���<.�n��d<����?���&.��hG��!�k܅�1�/Eҿc�<ۨT!�t �]�e��q��d����c%g[��s��;����j3��\$�B}���h�#�b��8����8��*�l$3�3�a����l����x)V��i�/�S�jb�2�﯏��D�%�yp�����"��.N��L�]2�b�v����Iha�Yer�~PY������
m��[�g|8�q�\g��g{��-���aVx�2��s�َ�Wؽ���(s��x��O�d)<%�mj3��PĐ�ܬ!@73+x���U�e6o��鋑_�����\D+�P���㧥������9��FZ����)��:E�����q/l��V�X<N�a&@A�.��4���N�GR�y&�E%���ta�p������j�h0�5��K�J*���_Vi+\�kK����i�:dt��b9��cr3Ò�1���&h�A����P/���$qpp��g��ܦ��Y�,�rO}�ع�(ɪ��8'���3�0�;IVo�r�;�6��kl�c5vr��9��th�匞u��w4��M�nl�m,b�,�����bL�+�j�?E�[n ==�!��M�v�-���M��E���PΠ�	��ᡌ��-��m:�������
�<\�kbG�sƠ���r��#�>Xׁ�3}\�3x~S8�%��ȨMkӶ�J���WI�?6�-ot��Z������h#��aƗ�6��s�A�8��]�i��M��91���d{�d�~�]��N>��Ơ�w�.n�.Wx�F�\��eŹc�6f;(�u.}��fr�����y���Ǉ-�Ij`���a~�ݨ�
O�h��q�VbC�QO���2V����?��b���uRTpC��������C�\���NaB W�r��{*����ꃠ��c=��c;���Ѡ��J���[�Z�xV���JԼ�l�3��F�X�?v�"�:6�iD�r�r�8��g���#��`'�N���W$��.��dly9[-;<�]To�O��T����4���xװdP�͖	^��э�������!�v�[�w���q��h�N'���:�Y4���	����}��n[l7{=w�����xuH�'��w�T)�X�=��@��9Gp�Lt����R�yq�h`�
ѯ��_e�N�ջ�pM�D\*`W-;�ȇ����N��9�M�c.�aϣRS�ϡ��k���<-�ה��.߾ѵ4������>mKk�(3�6:�\k�P@����7>"�Z&FF5ˇEc����Db7��!��-�JUb��ޠK��UQ����"�J�ّ����au)Wњ���9<|��G��zS�O:�0ؾ��\�]��7<\��7�2���T`�w�����	C�tN�S\���Q}ی�	YԺU�������+7�;y��[�_�l�\�������N�b{i�IR��(�R�7��A>���$1�@��x�?�S��'6�/E�8���no�2خB0��1���	��5�@��H&���Nt*u���Z��(�Mq�q�������������������&��_$/L���&u�0�Z7����N䥏R��@��ՇL咅�%��*�zc�>��I��F�Cj�8)NS��^����g����o&�
윜�Q�)sn#��'H��e�)�!����܌���gf#�ߴ�����H˭d@�u/^�o����=�Hodn����J�ٞ\&3��D�\i�)�oȧa⭨w��y�J��𡾻$y�X���^٬J���e�vn������2�"�q�fp���展��ľw�VV��-Y-���ʌ|��+x���ۗ�{Xzf����LQ��8�0�8*��0����M�\�w��k7�(陱@�0�7���\��Q.�콁o_�Yc1�I�u�c����9!��
yrxg����_����6s�ܕKB=�DI��P#V-`�8	��^��^H���m(r�,Ѭj�~+S���4
C��2��O�qq�R�J���hb̓k۟Cأ����(Q��&j��wz�Xw 4�y���{��~<����V�_��'���=��=��76>\?w<�%ÕB�Ve��n���+a���u����0�����zt}ON�3�E{
��A������0��n�SP�%�4����#~�>|"����S��Ȣ�K�H��e&��x��<T�;���6���^.sE��{�����o�IgZ�Fe�9���Ǐ{I��ӡJq-~lq���5!J~~,d���#��w�P�%_��H�s՜c#y^��٭�^mg�BD�s�����
W�!�{�	 M��#�H���99��Va`�d�] �g���I���{_�c�"���¾��~Y�'��v��K{��2ē�E�6�i�ԡR�=ȥqI5��sĢ�DX�W�8���}�>���N,aQZ\��b���Y�Q���2j�>�k�#e��A{��ʅQ�Q���3Wz�=�o�q���T�+�dC3�Հ�=�lo� $��4�a���L�����Z�*��/���]EfO�ٚ/Yי5�.�G�ֱ3׆�>��iw�f�!�-ix�&�Poĺ���=����Ǯ1�����Y-��:�@���;�"AP ��|� �zK��)�9�T���Ů�@�q���,�@�!�XONN��%�qs��(�u�q���v[��]����%p[� 2�[�P��l)��W���>����Y�
�����X�}�������{���x�M:�.�{��0�k�������!I��ye|��z�υ"S�o1��jFVO+c!zs"A	�1U<�������2lk���^�bx����|3!��"N�X����ӑ�c���C۸����7��n�6�}����u��ۣy,�M�D��� �|����2���{pY+����a�K�މ�����J����eH|���̘5����S������.�ۙ�'�����w�ل�2�9Z�-�?��_C��/v��"y���}
Wt�r������Y>�B?ZE���N��6�߆+������h���@�������U���f�WpP�[��qW���<�zzѹ���*�&��=��MƂ4	��Ўj	.�� G�@/��Kq�����{mm�Wi�93�IOr<�^���$4z׀��%�eȀ��W7�����v�nѶܒ�JL{�w!�M���@{�5}v�=���'d�!&��������I��QS�ɽ���;%t�?�!Kp�ŉ�_����/]H###s��Bl'�M��ൿ�\��2�j����c/#��)01Մ�N�ez�iew����Z��Z�}�c]7�>F��[N��8��c_$D�]�4�` Hv������r�Oل{D
�XET�^ɹ�X�P�E�ON"� "��}�N����q%Hͮ�%uR�h����}�?�B��H����s������ ٕ�+��Pԫ{��~/ �E/�.9��w	�G[�����`��A�����x���O������-�&�A3������Z���cd��7�zw�VosG�9ϒ6]��"��`<���2ƭ^����K��Hnڲx�p�� ����eIDY�V>��UH_�8〲كy�5zy���ì��5@�D&@�.�6F�+�].>Kc��P3m�9_�����:Ccc��4������Äm&��|��zs������`Ҿq��7����:�w_Xgu�6��������}� ��)��ܬt�6|W��������A�e?���.�k�	�P����q_܅�46��� [|�	�T"����.F�-3������`�)2ݎ'���#��N"n�7���� �Ej]E��a��#y�9G�L������0��} �W>�1S�K6��c���;�כ9�9���@m���Q����j�� ..nT��x,�|j���W�U����M���j�]5_��nľ�f����i��v��? ��o[x�f^���ۊ%�6�ё���KŚ��@��7� ,�R��RTY3D�;vl4��Uk���@�80��qG�?��W�6�凭ƓT�]�V��D���@%A�|p���f�{	ix� a,�I(v������ u�5_��O�a����/pt�����C���\�8p�)�.S���R�9�G���#�x���~�\v��`C���o�j��iQ�S�\
p��9�e$�p�4ȷ��.hnoN3x��tFP��2����d�X�(��՗����߷`=�w�rOJ�����|l�g��{��!#vp�1�����v@�G�^ߙ4�?V�v����pʹӬٮ�Y�6�*&�= !ާu߻]�/�86��HEcY{n�F6�\�AԹc�>����H����f�s�<�k�sׯ%DP�o��E�:nzK�Noߒ�⦹V��@����v&�~>���:�!��vJ�\���_�Ʒ��U������P9ÿ�6�#G�Y�Ƀ�é�������$�����9t����-��6 ��2���|'�?ۧ^�lF��o�F�������ϷG��.�C��t$��R=�@S=��ǳ���U���]l<�,���8E̪p��B�v�0���_�P���d��Ւ]��:���V���s��hq�ue���k�LЋ��>�K�
5O-�-��?�A8�2�RFB$9�qG�ku��{�ճ���m!�������:��4�ש�ѥ_>R&�ef���P���P<i��ע�=<�<���v��˅U������f?��3�=���g�yT�Q�+��&�Ij���v�?Ɵ#�(�F%�q��e#��y���!l�i:��^"*g��$�ym_�����k�J�Ug���P�F/L�����ˀ +�;��������\yu�U�'�F+�� ��s����vU����ɷ�xQNt;��f��K.�\c�'uuHrS捯v&�Y9��:Et\<4>/*_?>��(�>����*���Ͽ��־�ߕ�	Y`�L��P�̆Ԅ��"Okhb�H$�V�|�|�(#�Q����{��{T�|BZU��3R6G�FʨBRD�yp�����Ь�x|�4�=t���S�י�4�,��'ޜq2j�Ρ��SXnX�,�Cp���RhZQI�1f&�2�c�2/�k[U��st1���[�2�\Jxf�u�[�P�kk.'eϥ&j�o�(Á��u����ڎ��?Oo�Tq���g3���M�C-rx�$۬��^� �87:�f���4�ng,��I�V&�A��9�N�sc2�T����@L�.�}��l+6�:�Pꩇ�f|�*;ҍ߄���2�l�K�,O�������5��rz�G�O�N���;$��qoX)�^�M\�9b �'>4i�Rje�ѿ�Pd:��Ch��Fr�������-�H
Eu�~�o��%�BC�+\%�A^fM_̌�mf���Sj��7ڷ��J���U��\�[�?��Z�
�6E��o�2��w��v��s����6F������~G��[�ї�z{ש�k�B|d	�i��P�RzHi����ysU��3�V�g���q+&U�WWѳsr�68��n���xh�čS��Ѿ;=�u`�>}��?�[�ݫ^l��}\����B��OŖ�N�=�~�;�@�
����$a?T�NQ���WR�w��ОZ�K`O��� lxj��QB�gv=��NQJ����3M��������.������{��&4?�Y�6ڻ9d�}�_�.$g�*�F�ˉ��N��"�=��L���K�]���A�V g����t,�F��[���NÕ[����ڛ#�9Pˤ��Ê%�7��N�i���yX%�N�Rԯ���;/�I�����UQ"�4���/M'��R"�y��l�+��K�8fʅ'妧�_@ ���7GGhw��%+Â%��cD��v�AV�ZeϏ��p����gu�T�+�3O��kQB�S�B́F��?�@-Kn���ՠҮ@R�f*iC0�ϑV�f�CĠ���������\���S[Z�;����_xf���+������&��.*e����ƶ�#���<���_�\kg�7J'���-��$��dG�A���r����^Y�р���p��va2GUM���z��&Mu����e�}5U�O��̶e�埌��Y�^i�jq\0͊h���p�^,*���bS4�7�G�H�[��ʿ��	�Sb,`f��{
<	����e���.���G;=���$:�L��e�L���[O���ҽL�
C�`���֕��I�ۧ��������>�_��KLۻ[�$|���k��������0$���c����OXc�bJ���x�A��qM�i�69؈Ӽ��2�W�����o��Y)��H;bR�#��=��Z����4H~>j"��8]Y� 'c��]�DB1z�F���|�L?��b�QB���{s(���n���E"!U5�L��6'��'[-�2���L��s����F�M.���J���`k镡��	�H�ȣV5�-t��H��O�|vM`՘��F�~b�Y��.A�^��ܣ��.|$Ŀ��V�WӋ5����~���!i���|�j���4��_��}�7r=�9�"���O�Kڸ�e�q+M}�$@@�(�>�<����/o\�N�0��}�n���̑�dg���usv:��>�+�2G�&<�?�O���/9Vŏ=��+_~�X|����\v@��_�m�nN3������K�=�p�a �H��bdS�%P@�'+py��d.��#)v!e��7/�l���������%s$⅋����н���Y��hv��:Ʊ+�e�#�Z?%��l�E~���9�g�/$��Sx��i��m�:7����hO)�|T̷�E���ڑ.y�h�P�5y�����'H����p-C���E�"
���Ǝ��uu�m�Eu�~eO��~NNJ�o�0����:1%�gY�����hhiۍ:�s��ֲ�&3�_�,:4��i����}*j懻7\~�>���☛s��7X~�zf8�x���W,yB�rv}��c	įnЏ`p�"1���>���Sm̝5��h	9�~~Z�>~��(�;�yR� ~VaA��8se��R�����U���I�Py�4��4�u$��1m�@�3�C�����<��U��}|?P�y��h�ۡ5�ƶ�W�S|z
����F��?�'��^�i񴤧ț	J��G�������5��B4�7w��¯�<9^�������z��!Xh4Wd�� ���F ET6_�n	�_av��s }�JO����^�%���z�Đ_�}-שn'����ܣĿUR��˷�iS���S�p���m��
�r~/h{�w��~k�㢐�q�V��`�}҄����Sᰔ'���5".}*��\�f$Ǎ���O��1���(�6� �}.o���������ϥU��;��̧��������V�N�2������8�c^�7��yS<W_������3��Q�ǫ{����ZJ�"�ݵWJD�f��s�}�h�n�x�������^+?jjA��C��z���Y�b�AL��r �f���������>�=b��Oq�[	'�<� �7���q���V�V��-#�̌���I��֘��`�r��=D�n���__�2}?՚�|�����eIc�'
 �ӜFLf;�P��K_=�\�j*��i:�x��^Vr&����Q#f;�%�N��_+m/�{=���;J��M�D�|J�\8	8R?K����؀&ko��{T�-Y�:�E���k/� �Rs�"J��QO��T�Ay���v�@aU`;�P����o�/E r���ed�%L�|��X���rX���bݝ����J��s#��\/���絎���げ+1�]�(�����w%�/�/��.�[M�l����TϧT�bO��"u��]�{��D'��z�XaRi�$�"���tHr�YV��)yC�t�q����"���(���T[MG-]!�ߕ�Y�ӂY5�������%��[��2�,�d�P��a]]�by�Y�-�G�?��X)M��eF�0���g�f~)�,�'���VeAz���'��}G,E�d?HX�oS���<G8�ocWW�56�����6����^���c�H6r�,J�sF��V��+��9^�9E����%�j.�����/�ւ�s?��8��FA˧c�s�{��`iɶ`��+��E�U]h����Ai�3bX��r� 4��J5{�m�*%�Q�JW6F�/L��#��WC;�NU�o�:�^3������@�a�.�e*fpⷾ���L�!�6�u�����\�8���6t���zN<�}BA�v�?
T���0�݂��[0y0�/p]�w�;::*�k�$�ű��i��k�n5wp�+2W�P��I�S��r��O	���1�Nϔ���J�mPTI���)�)�m�D��:�W2;Yz������g��Y!��\��g�v�i��M'�?Kg����qJ���8EER܋w)A�S���݋n��[�/ @����ڗ����n����;�gw�3��Us�l���_��g�K�E���	zm�s�k�q���A W�{�h��z�~��-ص����Tʏ�L\� Y�*�X��[��A�g��%�G\$���V�QB��G�U♭���f�\��#���=�'��\Z ���Կ���Rj/��{��?������Nu�."3�� �)�g���>R�eO|��w��@<"��]%��Ξ$��Zm�6���í���G���1����[< gW��y] y�⑇E{�l�8��:�sR�e�35�����l�-AWx�4^��Մc�`�+�d�g�r[��yG�'Lض#ӝ�FH�"�/����u�S�N��<+�L1��L�m*������֖�Q?��j���������-�KM��%��H/\��S�@��7#3�+�Pom�"�*�d �2���w?��.�a(��br��Qh@�>�6�%PT��?��}����`M�Y�B���S���Ѧ�;�~0�j$2��lL�	�l�+ш�D>Zm+�lu��'�G��������?�19�3���ܞ�׉�B��0S�zn�ˡOm�<�L���,FR�"c���X��dRjо$3ͷa%[��0a�ĝ:�UFf*�k��Ҩ�lr�S�)fX���}���|RŸ�4�v��l����'�������;�̜���Ic���-�fO�%	?~����:���]L�������G��ˁ��c�t5ꔥ�����b ���f?f�s7sT.,��o�Mj��$�띥��k����&!RP���"�N�2��7�_}��q�Y�N��\i�ؚ��YLZU
�(R��܍ƚ�`���V
�J�?�<XǮ�fd��\��1��Ye��_S���)�͡YLfO����jn�lC?Y#��N�ӻ�#!�;o�MSd��o�4��?b^g�%Ӭ���
�IX:�AM��d`�w�U�o�0��Dn�L�eX���0Q-= ���jd'YՙkN`��Ԇ4@K�"[n�p���X�56?5������:-x_����Q�����n'�"���1B�M|G'�-�h�^2��@��4=���1!C���W'E�;;
ˣ��cU\�;��IF�z��ѽ���N�_x0����ߧ������1�/"i ��z���u��&]s=>�����dh�M�����)��4eD�.���enFpMLjc-q������%�?�չ�v[�F��%�������D|�/N䶷bϚ�4mR)�3��yi���p������vQ�=7����:�}�/�U��<������ȉ�Dдg5U��<�h����4%+�����_%§� �h��h���g���r0t��E�ҩ
/^տ-���t��q䡒#��W��'	�����耻�o4��N��^5�vWn~�U�V�����q��Ο�Ǻo��<X��tt��[W�GG���܉�CO��/K��w4pAA=RF���	\y}[{zi�"a��/��F�H��wA�R$�+P~�����"&Cz�֎��a��-���d�����EE����j�bB�<�qLF���3Y6cx���ݵGtyVG�M�_��,�s�n���qf���Ϋ��	ۼ�S��:���^j��O�����L�{-fb�D������o.��Cn�Lu��]�6�e62��E��Dk��椧Y4Ey�It��+O�,62����$�80O��I��$�C�߰1`&5;��`�cmOAqk�6 5��vp�{���l����DU���gABHs��J�E�b�5���{�/e�W��ٻ"ҲRA<�]u��Hx���1��~"hR�W�P$ߪ�4�c���\�L>^�q��uwk`Ʉs8Q�Me�h�8����F�M���4���6I�?s�h`�gX���&d���O�x���C��1���C/4~��D����6M��V>%��c��Uգ.մ���iʤ�; ~3j�+�7�"�>���FE�ߎ��g��ĖO�����2�ٸ�)��Xc���>/�?��,T4����w�wyCf� ��ќ1!UJ��d�I�7a�M�<�.P96^��ߍ��7V�D�Oy����������q�5>d�y�F�,��.
�d��N9�ӫ&�q�_���Ye(�M��{�����F䬚�B�q�ˤ_���o��.:�rd*���J�PὍ����N�"Y��v�@�B04]Ρ$���P�:�f�X̐W��P8����x�XT��`��H�;Бk��n�_.W ��ץ���ȟ�	*f�~�5�!Tή䨣������a�y��N�����}�Ab�W��*V'���W$�L�/�Τ����>�s�;Ҋ�p�!��ҾDT73��̩��`�M*9s
�n��M�� G���d?� � �9��~��8
����2�7����_��m��Upp�w�i�)%�����[�r҅:�YD�sqc=�w�,�b,_�1Jd������nҌ���ɇ�I��C���H>����*�7+7^��ѿ����WVW��!Q�_�Ro��7a���Q��$W�.��M%Bwrl}�����x�/���[�b�����Fa�|ʏ�1����~���K��PKe�Y��|���i(qۢwn��^��0�E���Th�ȍ.�kPH�!�����;��ז�(c~�*J�r&���I 2%��;	Uݝ�ܵmx2,��/p��ҫ) )���fOSD�d)׸F�qG�q�1��N{�+�Y�7-	,��i�Ot��p���5�-��}XXDaV�9�,�t����BĿ((RYz�?`=���~�I���3-(�c��RJ�#��G�3ޒ#���2����u*q�Hg�	q�Q���'�}�o@b��a�~^����Udc{��N(�k�|?�ӼӍ��9�{s�ʆ}��0���{��r�Zx��Ү�T�wy
��X�LЯ!;��C����կ���JI��8\"�^x���#av����.��V��ɩ(�Z���
E�%�7j��GO� Q`�1�q"�`��0���y������;�P�?7��֜�~uZ"��������.����vZ)��w�[�K'7"~�I"S��4�����w��x�"�t���ndK&A%�}/[o�d���A�p�Ɍ;H�&����k䇮�3����D�B��O_��������Nu'������;�Ծv��5s�/䍨9৩T`@Į���Ԩ�ZPQ��\:^�<,-G����<�v~��5�b���ꜼeU�{����� �π�q
�+����&Gy��X�mʪ0`Xl9��;I�����T~A� �u:�fBC�#����)<~����OZ�����@��#+�{{l�Ӻ둤��jFg�7h�t��p�.B�$s!�_��J�OA��,8i�}/��|?�ĥ�Xc�vpv������1[��⛈R��%���c��g�OW��X�5%�6�{;���LAc�����a��`�����9��ȷ��Z�%#~+�/O��c�RGhd����A���U��RȤ7�=7�����m%�<J8N�9���5�Z����v;]x��P��#9�9:L���\��(���/eպ�� i��`zi��|B���Q^�����5�O/���C@'\ڵn��B1���Ϟ��'{K�Q� �s��*��j��T��~�}~���7Y��!ԡJ8mR�4�^E���z��f���MYh��� O� _e��Vӂ8�`�M�c�a��A��&�x��u*�}V�z���s!��7�YQ�sq��8=ȃp.Jy���Lڌ!Iא1j�7�J�&&��@���hw-�飠N�e_~��?����%4��舢��.�7�`Ka��v��/��Hك�������m�Q���>�KL��n�a�/]Q�D�Irj�q�(�c|�2���I�o��c�LT�8|P]yd��%߼�ѝS�J+�c���,��ݽ+cW>�Rw>ZYY�|ya�xP΀�t=�7�/Mӊ�BS\�9̢�m��W��>�n�^�m���~���3���f�Kf�QɅWUUU���޽$���W���Ͻ��� F��I�nR�ᎎ�=�;��9P˖7-g>L?���y��b濆�xs��s�̳:��^��,���k،�#k6�M�?��z;{�u5i��n>�l$I�ݍ9��^�@S��M��mRC0�s��ac�^M�F��x�Z�i�1����=O���s
i���Θ膔�E�@RXIv�fM=:��\�������>�gT1����/�zj�-?B��"n�`��/�,�űf/���5���7��g��p8�~s�}����$Ǐ�o�[�<��erl�Tԧvk�n��{oiA��̰���uNl�y��D��L�H$=���%���Uy�ajY��DD��=��4kV)A�����R�Ɲ�ZD���Gk���;�Jhe������V�[uXb�S����
�t�W�Z�d9»YxF{��x&~��f�ג��$6�O�mj%p�ϴ���y��
��f�U޾עV���8�E8�����|
��)JP2���u���W7ț��?_�����R��g���2�	kH
ʳ��6q$Ͳ�q�p�sAW�x�q1Q&�1cQ홵"�ٳV�=��L�SS�Ͼ�r�I	���!�̩�X����,��0I���j];��������е��f&w�1/V���'�_���?_
]�U���Bb�稭�3�j�?y�UJ1�뗗i�>l1^ڻ^�A;��ь�� z��$fUav��-N {���z��%�W�����:&Z���x��C�����[���I��,�a~�l��M� �k�rhU�է�	�7��xsU��UޫwB���jk�M�X+� <��+ȏ^|�5H�Gޘx�#GX��$0��W�2����J5:�ef���6������0�Ͱԅ<�>ݬ=<�{�k���b>��M��.�"�{g���0��q����ފ�N]x=�󏰌p輏�/x~����W;��[F�s�M���vi��W�A�;#���)@���0ߛ�vQ�ܖnzM��z���/?̦3��.��ԝ��G�=�B�d�z��A��?�Gi\K�2Z6���|NP
�m��֗r{�W��f�e��������x8X�����T�l֦k��w�����#`��Ǚd�;�!�.�)��/=�.>.�.-f�+.'��LU,���:���|���w$v/u��2�ui��U7�E�'����/��ʆ�S_J�.(��|Ϯ�Hj`����Jj@�*�l
�H�ݐ����RK��
)}�ճ>ޤ�v������&=����͚ύ>��Tw�oG�_]�%�-_�]ǻ�J��v=�<X`W�{��ju�lg�tSΙ}�"�,�k*W͞���� =����3�Կ��P�1�^6M&��_���Va�	=�ZBw_�>��_��\8hY��U8���Nl^Q/���VBR�	�����	��ΜL��?#q9a�Z�����w���\JАg*�T�\�dੜ��aT��RR]�?u4�I��tG5����u�FԧV�N1DC{ܷM��ft6c*��,rq���EpF���=F �"���vN(�yA����I�䞯[����E�9��Y�?ÓN�9b��W~�.���m�<#,�o�hdbC�!�w����۷쉯.��Z�e�d?/���bB���̢�6M:}]���w�vo����j�6��D��J�6�/�T���333�jǗ��
�W/��g\�U�&D��$G/l�qwߢ��@Q᭧�խTU񲺘BǕ�H�Ad[L���đ��x���TԴm&S7l�y1��b�dG|D��CV���zZ�~�9}z���_��o�g��B���vp�����y�0샣#�G��'�$��X{TiQJ�,��M��!�Ell_���P�#����u�ތ��1�����"oc{ٰ���5�:x�!�g-��(�Y��+�2�/Z/�s�"T�j���_�Ť�A����S1k78?퓮���zJM����(QC���ɫh06G4�|��^�]WW��^笥PĻ�6@~��nO50���߿�s�G��QCf�)���D�o�^dǝk�<0_������<z�I�'N{{�=V�ƽb��K���-�8t��3��м����_A����y�kP�cKM��Nzx��4Z��7Q8��gE����M��y�L���\�V���iqP*�ۻ��L5¨�S�8��֥q�q�9��LԄ��[���E+�a��MD��^GX�n����@�u�G'�8������u�aʑ��7��;�쇒�_��m�1^bd�|M0�Q�W���iX����/��`�U|�����1��E�g��f��|Jy�>�gr7�@~Y��&f@GWb����gNURJ�_KGs�E�0���l�/ڷ��X�7�U�N��[Z����_T�5 �qL@�i��^����J��G�:�Bt�@����	�����i���<�|����������$�.d�tcX�\�o�5	�s��J���i�o	��Sj��d*vb+�����R���Ծ�c�$���﫦I�؎��#s�ߩ緅~�ѿ�Ub}�2o'�E��)��R�V���J��y���M��9�wȿ�Ac�[Y��_� �f�BB�O5��24��`&���5��<��ڍ,OO43�ϲ�����q=h��/h`@�����!6y?�%D��@-&<T�\��3CF��_~<w����s~���O=�q����$�U��<[�{���+>{��z��WLu[c{�'��+�����v�[)%�W��N�
���f0G>q|slIo��3�}k7�h��F2e����Ճ?�Iן�͐����j�]�x����Kg_�*�k��5����ɪeY�p�O�rԖhݗ�?����_�����|&~�f���2�����sxr~����I�#;È2�Rm�&��>�����Y)X؂�Q�C�V�qjCX]�=�#[�J�6}b �Ӈ/������Ca����?r��\�/K�Y�Ϥ��>�&��{}�����4=*��q_�6���C��l��ܥ�dk:~�>��Q�9�`j!�o��b�~��DG�Y{�����,��mv	������"x��+P��V�.DBzuWR�fV
���̭r��H����k��Hz	]��*�!�Q����x�'0��Wb�����ٷ�����6���z���hvߘ��l뉴�>(��!��v'լ���^�!]�_�*�BN��@E�eU���^�NQ��> �h?�Ҍ�%3dPTI��Ȍ#��;r�Jp������p��Jc��>0 '��z�ā����{�\�|�4����ǒ3s��J�ƕ|1C����%���*������>
��x��n�vj�)*�|sMxm���S@�e[m�L��%��G����¾0��L=����tk�����>S���(@4��AB�`�B�w������ʸ�Ȧi@��
W�i��'�(��Z�N'ĩ�����)����n���-kУS���)�0���;��up`��u'������ui���D��
HJc�U�yM�{P�������ޫܫքEs�a�`4@ ���}����� ��SW��ڃ�Z��*-�B��r�v�����E6�']O�uږw]g����������_���"�~c!������/��7/M�,m�Lr����*�S"����`���ė����Z�����L������t��b795}�K��������o¥a{e$qɾ�^�P��&G#���x�J�����C{�'������o��wޘ,������x9�V�Q]��3$��VxkF�@�x;��g
0mE���U���d��Y��UB�"�2��a�._��<�t�pSF�zt����R�bK��l���jk�\��k�m��i]j��T��jL��y�ZH-˔+G�M���j�f�`��h�E.��#/��!ɗtL�x�z�������������HW��s����;m_��I;*����$�Ѻ��YI��.��PZ�ks)ƛ��?�]�� U�s��Rް�	����	�sH�4���W�b1f��&nHYb�kƳJ��:�����}07����i�����C���Z�ϪS��v-�I3��X$N���*O '&P��pK}`1�3����
Y��Q����o�R2�l����k�X*�Rv;Q��f�oj�IHy%�L�߇B`����{���T;���P�.�Ύ�ٜ�V����X�*3��ж�El�>P�����Cry#�����uK,�C�=�<�ö7��,m��m]ԡ�N)�o�s��!�*s��D���1V�V�8�Z�b�_�c����?k�����ޓ^"C�)|C·�5F�ݑ%%�		x�]]��ټ�fU����s:�m�޳̽�w��-lP��Y6�N\6��ԡ�x�t�!���	מ��HڿVk�ׅw� =Je���_�݄j
v�F_�?P�&c��}w�����r������S�W�rt���ĥ��lOd�Rh���`�]>��̼�=��Z����3�R����k�2��+��$T�\-ܮgs�I�Mď��hM��_�о �G�@:�Ɏ��T��+++`��Sl�߼߶іK)����L.T'��n��HMz|�ۄ�ǠZ���7�b�3��nB[CdY�!{f�bR���N��zk��2��ca�.q͟üm&��vBl��ۄ��w���z&r�9.��;'t�T�,��ľƵ>���H,[#o�X�SC�U��^5���9ޘ�Ni8��6x�Ӊ��k�O��ǒ�[�fyrd��W����P-���	Ԗ��1G�4�R�5?9NV��\���'�i�S�C�����	,C�l��c����SNn�P{�b�+�ˎY���h0m��ĺwLM�{i��.AG�����5LQ���a�\�/��r���y���S��ėJ�flC!TE6�^Ō:����W��Q���x����k��bӐ�C��"�4hMvl#�H��ҠB�l`~A)m�.��5:eJa��z�[1o�{cA����:���4 ѓ��a#c��Y˨W�Aǡ����	���4�9RG-�\����q^n�A�e�?\��O����i��48\y�ߋ{�-PԸĴ����{��w·� s�Hё�6�B
t�3��c�u4�W�̳�nś���_�)S�U0b�E��e�U��Jx��¦p+�:��<�O*{��0��'���3�I��>jR��W��DP�x�V���o��� wJ����Ŕ����˯��gs�ܫG��R~�>#!��ˍ�M\������?x9ޟ�u�u1��q4�t-El��\bl|��0�乸�l=�M'Y���)�l8��V> �Gm"��Gw4$�SG��{QN�nhr'"t�v↥��x���`S�0������VT���ߋ�w7e3�<�����!�=�J#M&������b&�-��|آ$��$�S]ib ��&��h��ubP.��w��9�y��'��R���ކq(���Vo>��M��H��ή�C����σP�2���Џ%�F��$�����.��|e��)���J_=a��5AЈ�õ�썶��v�or�ґ�Wm�R������*����>�k%XDӠ�o��HS���H�`YE�#�p�N�[�n�P�h.�a�wt��J�ıe�E��&>�1\�+�0�[��Eo�����qU�&Sޜ��Ȫ�-�T���+ּڽN~
���}��x�*�^�?��S���f�����JV���ıpND#�{�cj�.!.�|��e~!tN��b�W�9�������&Q��"0h�q]NNq�%gΰ��:���P�0���V�#��=vRG�t5P|�����J���{3���=o<��(���Eʰ2�Ώ��Ȗ��'�1q�?G���@�K�)�S���)t��1ʯn����	D`Xt��R�B�+�3��!���8��{����9�ON�n)i�W~�}�Uk����>^&EpN��ExqO;�+QN���ڣ�<��ZW`��%v���hD(�wN2�ۄ�F�o/9�\��d�ƚh�������ҿ@B|p� ��`@mb�� �̰h;Ϫ�>�����߰�`�.��Ӱ
�q/j�����)c�,_�F�ǵ�϶��-&��N�l��P�Z�����w�0���-�H�k�@�⬆]?����y����=sO��\�;��^��Y��! ��\��g�/�
9��1<�Kgb�^����4�"�
k����@.���w�u�h����Ia#�?� ���{�4d;;s*�5x�K�a��_h�UBw���D��e~�w;���.ޒeF���j�4;�ȥ�ȫ��+��M}��R�-���n^L�o�;}��(�<^�� �7��Eĵ����}��`<�m*��j��kpx[��wG8 �R��v,	���M���q�X�l��� q���7�Q�V^i�;�>lM���Z��@I{��;R�{�� no�AĒ}¯�b�@�\�]�뚎[�Qvב���ȝ�4/%tP�c��
k����7�Ӂ1��+�Tn�M��1L�o�%�ԍѣmqcMmx�i���zF��6��×���	���r4��8����b�L�	��h�1�O9�^(�?�=|ҭ��)X����9��!`����zh����o��"�`���#h��p�� d�F�*��G��ѱ����"��A����s���]�+�ՐIG.:5�l��%ߣ�牋ǂ: �6Tm�SB(���[�]�	���('W]��j.����c#����p\��i$�0&�~�V�u��D��'Q�FAk$P֏E�\}F)yH|�K�(��?��m �gѺO6�i��%��c�>�|�����v!Eؼ��S����P��%���5;k�ϲ�v���[��t�C������LF�.@����W�Na���caa��_ �O�$�ݚ�*��I���m*�HC^��n�A�V/��z�;��� c���^�E���"�$Ĕ���W�E5��2E����������m��o=�l���@g*)�OA䏟4�H����}H2�(�AOAO��8g���_b����o��'��	���q%�k�o&=}�����M���ɸM��Ho�&|§��Y��7���<j�uV����r�O�������N����2�hS��bU��!���[l�Rio��b��K[,�%�湷�Sk��!O�_P#�CY�a�)��NӑI��ָם]:_�B���I���>�G���E"�"^�H΄ ޷�<��`|	�C{\�l<�R�1me =�[zu)�0"J��`o�+������J�'ϻ����,��1�Q?�[gg���
�g��0�aq%�� �����ɑڮ8��v����:��k�:
�{�z�A�fݣ!(����;�`�l�5���{�D���?�SSj�֝DL;� �,t�i�J|�h��䔭�2��zjL�<��zc2Y}�FK�7<э�tm��q��gBP9�9�0B���8%ǧO�*<p��U^�Ț��P�P���UW���P�\L�yl1J����k�I�\;�FnnnR�E�������q���s�v p4i����iq���8s �
aW2)�����m%�]�]�5�Ϭ1�rk}�E�Cw]�k�i��.Z�ק �O�Y1h�ͩS�1�������9	Dc倢���	�][�����"0�h�����U]g���bFI�����{7��1H�0A��sz�6��u��3��;p-(�X2e�2=fމvM0�S�Q$A�r%/���x4��X�����Z i8�qE�bCx��2}��N5��5�4F�h�UP���g��{�����Sy�{�u�u���w/�ۘ.�ڏ��.dhx��鑪P�%I(�����P���(}#G"/���/�-G�!Ce�5��'��]l,�M��:ӗ�,��	�$�J|���E���:�-gv4)�ږ q�1�U�*�*6.n�Ff-^�bV�moI�&�O)�QR1;GTx�I��U�������)����!%��8��y��4}���!�ɴh۝�G��DyUI�\o·/v��&\�������?,kw�ߞ�f,�y��������sW�^�vP8͞�����t4�0d?y�� E�$ ('��Qc,�#B�s�Rܻ�]&�I}��w��HMK�D-����#C�c �r��q3ͽ_�dɇۼN�j��3,��P����a����$*at������B��@֪VP˓��xԍ/��f$�!Ƭ�6g��bBk$���W��,�g�t[P���chWq�������3�HL��;M���#4��*٫�讓��!{=��d`�qT ����1����R0!E[m�Ɯ�՟�N?Y�IBE@��>*��6Z�.z[vF6�i�'㤡��8��Bע��T]�C�A*���(q�R�m2\�2Ms�W�������^R������ʼ?Ǿ�u|����ZA�*>1!&�ԇ�歮z�"pΎ�j�/�Bp.��F�b>$�rT��<���[nuiگ�.@�cņ�j��厵�cZ,1��h5�	ͨeBI�2���+��3͜�}�H	�}�H�:n1�p��!��e7]�T��/t���G�������)�xȠ�{�쬭�z�
Yݪ1��&����⬖H��A�DS��u�:��F�������G�d��RK������ԭ
�#m�*��}H�͊�y�W�6�n�hBrH���_O�⒇N�M�+�l�Fk]�wԾ��Hz\�'|�}���zML*�����A���l��{�Y�0`[(1�V�eW����S�i�K�0�mH����}�'��� ��$P�Ċ(9����Z�p-���l�����w����޷�%;C`��݂;�Թ�$�o�B1��H��߯��;�����v����U�>&҈<~�7��>ܝx<�zLKɋ�����h�h,B��$8����i�x�B�wJ��,�J��!�H@�E#�4%��*r ygg�Ba��������u����{􆵌7�V����cl�s���D��@P�_JYȥ��	�y#�ۇ+"�����W�*�B�Z 2���!�VV}csS��s�/ P� �m4v���;8 �����W|��l
꩜M{}�F�?/P�6�+f|4��Q���Ǖ�_(l^�n>�ٟ�aZ���>P%��MF�s�HЍ~�-H4�b+���وB� ��z���I��
��Q<�!VV��tOkB�$@�u��W���[2Jy�q�j|��
��֎Ѷu%�>v�0g���:W?�E�����-Vo<h[>��d�%�l�����$=<��{��d�@}sY���`J�4闚&A�1�/�fL�i��2�z�\�7hV�{(tc)4�Ƒ/�S<h-c�#����ck�A�Y�'��Z���O�ǆ~g0�����&���[Las����,j��v�3��	�9����&lv������"wcfs#��$,�٢�TJ�k�~��9ULG������Q"+�tm��Oi���ŗ�P��9�RH��A�à3J3���Ì�yj�S��]��*z�t���Wy
�T�l�B�r@��/���m�O�@���2�T	�L�B��׈K����3k�CI~���Y�|lI�?oX�z^������%Z����MV,#�@Pg��K�(GԻ��G�h�tv�Qdf$k�����5�}������t�j��)@IM��Ok6�]����6�\�u��Y�y.}��
b�6�Jf��
��u�~�L%�V�q��*�����ԣ
hןXTV�{�Q3�m� "DR~w�CN�8$?��Ε�����Iʾ�e���aȪ/JN��&5�e�}�(����us�����߾��-�3v�[5kj�6��o��R���x%����s���S�-�?X��%2��G��U#P�
����U�5�-099�NJr�#h�ޯUS���t*��o��H=_��������`k w�^�����ݒ���yT�{�AI��k'O(	
}���<� �E�	�|�Q��9�~g�rD�ŗ��%Q�=O*a��!ǋ������ ��m-/�榀��_���ա
f}�D,O.t0�wxmM����1�َ��%l�cN�
?Uf��IZ#�f������G1� ��ۯY�c�ʻO[<3�i�e%^L�qMM��cݭț��)	o�&�y�/e(
��$��V�&&	��e�l2��e;5Vl�m���k8�\ku)mr���,aQ��M���4�5�L�o�p�����a���t�6��ZǏ���.T��J}�>��Z��$��l�l�LF�8&�K^AA��(G����TEi5i˵�fS(_iNA�~'��̬�`i$��%L�:�4x���T�ǡHj<�V���������������2�s>|֓G���1�h(�#�u򐚟�����l��BY.yU���"%8��k�4BJh|�N�=j_t�d���1f5�fW�����ڰ��SS�ׁx������睸cs�~W�����a8��K�`v�␡1����`g�E?DdJ�u)l�<�Ü��>5��"N@��Yz���Ґ��S���D�$��3囗OE�ZV�H&���K`���-�^����2�[R0gͶ!{˵��aU4�[k[#��j��O�L���I7Z����j�R|cG��gXOo�m��?-V/�<�:��Ȱ$����3�Ѷs% ���f������U��#B�Ҟ8�Վ }L����V"���,0Od��ʷ��{�ZDʄ�u����%����J����N��O#oy��xe�uNC�,e;�`�3����)C���_�Έ��>����Df)��i�J����w�5k����HPY������dF��+����qݺ$��_/���~���ٝ$�ʠ�N.�A'>��$��f�R���3$�s�R��2��%��#���*����5[�ak��L4a�<u��?��we�������Y��e��� �*�o)��z�G����R�4h��F�#K�`"�(�x�_�b+��n�ŀ�я����0����V���wzW(|��ahDnE�����:�L��2�h5"$cp`A�h��D�1h�ﳫ��� Z<̗�gz7�s^~��ϗ�1�6Ww���B9_���oE c4Ƶ���cO'��W���y�d'\�-�B��8�B!��+��0�B`���sc��֕6ˤ�j׊$c7���X�q�e�����<��0(�_ދ&���Kْ�|��D-��9�Q��2�W��aspG?ݓи䑦��gȨF}A��ֿ�IFP�'a�T��'��*D�� e�#CH&yF`�fr5�����D�z@�@O�a� �M/���?��@m��읶8�R�k�8K�cK R:U,J	���=EU����A*ִS���Y��Ӈ��Iw{v��m�����{(�
V�fy��� �Nl�wqfiڸ�6��Ay��@�k ��!�C&�l�-�2m�׹��)�,+7@ӈf�S`�oE��d�=ج��URLs�oH~V��"ك?����5ͻ�������=�Imp�������4�ɚ���iX�O���|	�MVIm����k,�����k_{��9!E�n~��"��!�2L��֔7�@A?�����pt>yF'��̚����6!���X��Jj�t����:�>�=<�m� �a���[��)թ�¿�'O���K�Sӛ�q�L��ޗQO#��77� I��Ja!nD_J�kg�R�gS�S��	���5]k�w��{℣1�?���4��h#+�	�vp�?��>~$�"cSm"x;Ω��X r���
�gթ�Ԑ_W�7�� |k7�w;����j ;(��u?9�{=��?!�=]j>{�(.��2ݦ��:�D`0`�҇����QA�����LD���C;�
 q�@HεO�̒7{3��Ҵ�ԝ��R�i�y�W:�
���>����m��µ<&7J��l��Ə��� �`�_;�A��G��E��	�8�c�uN����ӝ&:��{'`o��C}��
��* �㘢}���G�����s�L�h;�XeH���tF�^���K�.Z�j.Yb�ǀ�x�BQ��(~��t�m[���[�b�c-�tUT��<����F�@�i�QԈ٥K1C�"Q� r=p8Q(�>	k. �l�eP�-�p s�Q����z�5(�˻3����m��T|�P��N���u!ܟJ�<���"05 �����+����d�D�!�J+ӯ�6{f�j�'	���p���B˶��G�Q�l��|* ��F�O1�j�N`Τ��?�А�asi@�/�<W��"���7�<���ǤiO��A�����k�M`&z�/��~�浞�s=(��
�
^��-���të�K���������MnO�jt����k��8ݝ&!���Fww�A$%�A���0Rb =&����@ҏ��o^����N������;{�9��_^Z~G����4�$e.|Š�kW���<DCm��t�F�/��]����Y�J$�ǵoc�͔F��'C��z�qR�b]!`�~M�%�l0�d�?�\�G�E���{���CDLP6�5'��Ũp^�V�n.�����S ���m[��{��~����߿/F�9���ȝ6���-�)p�&��i%@�#��=~��8�( �5(=r����i�;�e�z�Ю��"�P�v>N�XW���f�5��)˫OV�"�1��1ܤk�~�2r�kD:M���K�Si��]�wr�Q����?A:�v�j�"���_���r���Sna������V׹drd��~�-ֶ��	
s����5G�T���\��49I�>�ݕbLO���b��/��a�hw�u.��g�7�K��(f:s�2�{�oE#"�kb�������i1�t��w7��������Զ��DM�5{T��cT�O��9!! ���� �����-���J(U��M<�F�M�F7���� �#�\^u�ꔐUؕ���ؓ���q�5o=�߃Cn嘡i�I�g=�*Q��8(B��"�S��#�t�/�w��fw���T�l���@��{���#iOY2�QQ(�;�;L�Դ`�R��/3���k@גk�;i�ڜhN$án�t���7Ө�Y�ͥ$�	/<�\���H�U1�� �&�(͎kg�;�V��v5�Ή�=-t��ڪV�O���թ6�7��H�]� ��D��]M�%MJ+�O��\��u 	ƾ�`%���d�ȓ͋��u�Y<O���2�{��X<X!Z�_��Qq�٩q�xsL�m���Pq;�<�\�S	D��ג���(��ȣ^����_5�^7V���>��l�����r>01�ßυ��n)VM]����R1x���uΦ�D�ͷ�5�3����旽U��\�_�4��.����o��y����ƒ�X��aԦs��&Rd�L%�.�,����Av�9B����N,[��q:��3��J.��I{L+�^Sj����e�qԱ|����ۻS9���>2��c�����X\\�0|��4�.A!c����Un_L��~]��,z�Xc/��������h����5�3Q��޶�����֒��	�P�_�k����%�[=+����]�1Ut8S�sB��;�FD�g�b�%��ə���^(�e%l������bw3��2ޯ����)�Ⱦ�ѠՄ��sg��n�� \'
v�e��J�B<�4hI�������d���dn��_n�1�7�c�=r�\p2E�A�ͼ����<B���u��>��>N���Jgø�bu��W~�ٟU���L�xt*5�y[��XGVG�Jr�"}%�-�'�;��W^R��㌟D�za@���ޮ�9OA]���q��۷�K��"�l�7�U0�9��\7]��)d^P�2�45HP�`�c�N��Ի�`� �5W��n���3��d̺�j�v%& ���8@�q,K>ٞ�`�x�����dρ��$�!=��>Mf+�&�Ё�/�Q�w�w�B�'�e�M_~c�XV�kpS����b՛�%�]"�ʛ4��?�N���&U�3rw/�`O�ʋ�7�	~]��Ct�+�jՍ�
�N1�O\�%b+rVT;׏rK����&�I�Dϧ�H�]�2�$%ۮ}J�sA�E>���<K��ʵ3UiG�O_	�oH�*b�~�&"lk�ZAA� N�^�Kn�c=[�ą��&���z�bc��ÿE�%�w��,|%S݊a���'��tq�644u�9��-�J��*��|jE�n?s�9����O�ؚ��I�=�?n��;�_srO����2hw�z�Y�Ej)������i�k�(�w���a�OY��|��Ε���{�����͠�?�y^F���E�?���t�4,���3�);g��˷����k�^n,��T�ӱ+{W�E�ޱ�PJ7����nE��.c���GW���Ʀw��<:	�1���\]X��d����.�=i�ӧ%`~
�=�%3�i.i?�7}ɥ~uLU%�)��Y����G�	�����h֖�	R��yv�(�R`&�,'W3Ħa��L��Vx�[֥�����n���⩪'�n��H6L��zZNQ^K�]`�%��z9#�7���~ޛ�o,���+V( �m�P(_�`t�"o%���y��Q&����_��˼�^��WN^9��in�Q¬��h֘�Q$ϙ��
�g̦߳cX��[?)���x9�L2,1�����F���9]���`otv��O�k�������Xg.� y�LQ|�JE.l!�iW��ϼ����א���A�s1���P��`�;0�*;���w��� ���w�~/��� �{�}�v:��yh�
0�V|����w0?�y�����;]^w˗!-F�ŃW� X3Y�I~�`�Dn��(�Q-�tɖ�]���)���@J��i^Q���w���k� �������Y��l�Ҳd��	�:��u���yH��P��i;.�R�q�Y{�J�����q��:��I�#nB�?��%��O����fkM��R��AG{�X�I}����a �¡�Z��ئB�@Cǫ޶�5A:�t�	\S�[f�"[� �kK�U/���;j�Vw1@�Z����[gEc��h4�c��e��T8ftر���rq�{r��3�m����"�Qy2�L�_�/ls녏�f2`^w ���F86���Z�@��� ��^W��-�;*1�>��A�v�uwW4b�k����۪��us>����6�oĿ�]�w�3ntwQ#7��c�ˎ�?�F�ú8Jv�����7T>)\J��;w�Ҩ�x�ܬ��Q��	}�����&����Q����J��k�+����#�J�t6�t[\!ƴ��a�|(�z�*DD���4є5����b�/Ĝ��-�\R�}��rl���3��ܞ[�ku���+K�������[!ȗ�ݠ���L"��ߢ,��eT�i��uo��dQ�~�l�jPd]����h�-g��E�>wW�ߊ����׷�̑<�F��O����Ȕ�
��L����;�ۂg�����y��9^�����Bӿ��M�H�#�ҥ;8㐔&m�}\��"�x�m�M*A��E/k|ڏ�8�h�,�u���uo[fM�/\�!���a���
�/�CѠV_���2OO����F��!�8ٱ��g��Kp�7��dT�c�a�������)������\p�bGW�	������4�t�����3�3�W����Dw�WJZWo���"�o_F���8��_�\�J4��ȂpW:�!v{3"�ꤲ�wM=L���g��UF��Zfx��E��	�,p^��)�X(�ٶ��72$��@���e�n�|d�H���	S���M�b��O��L0����p|�In:q]�\�w�%���q\B���ȣ#�����́fq�T��x͠M�`5��y�~#vcK骐3� �
����f���`-V� ,<WF�q%��l�K�ͫ��M�Zmb��PAP9KPS�k�܉ܓ��ED�*xX��\���Qakn`��g���C�J���,��1[�|�irw]�X���X1c<�F��ʽ�rU���ԧ��2��y��o�����ݡF7��U˲G��$�ww�6�:�;}��8+�(��ҹ`ob ^$UDl��� -�/?<d�ټ%�6*[g��;+B�8�2�MU���L��5�'�m��"�9�<!�%� f�y�ĵ�f�4�=��Լ��wzܞ������Z��CB�pJ�E���k)��h�<�{z��������H���g�E�5<R�Wr�	'���û/y�h3ZA*y���:����͌��T��`�I�����[��>��A���9�_p#5�o�W�M\T�z�I�<D?���gNS�^���_��$}Ei5R8:{��2^
e�_Hꭂm���ږi�
�T#�9����+x|��(�WXQI�9@s��2^x�)<$l�'A9"��F%"7Cn�nn����֊۪q[k���ʠL#V�f|6�'$�Z��q/ ��L(����V���$:�_�ΠoW��]�VF5�(�Qs&�
�?�����{4�� �0��ʞ�z�1,~�
1���"qk6�X���O0Y)7<:�Z� ����c���񵝃����ԉ.�c�𓎴]��3UeM���౭cv����0,��M�|�Z��U����pGծ[F	�k�(�ӄ>�м���p���+S�7ޒw,RM�x�r"/��DwTW_?"l`4������>�UX����Q999͛kb��z�d(�ie�\l��g�z�2��|V���j"Xٿe�i���\t�ҡ(�)��/�	�(��	P��Xu�D<�������K�in�ɥ�-3@����0�ޓ�ӓ�C8m������U0\sg[:?���m�� ��O��+鑳{N�(��@��������e�����x�H;�B������������_&oz%t�2�b�M3�
�w��)´��ɬ{lD���������N�j-���R*s!<���6��!���e�+��c��PS"&��Z���*��������_v=�g/o���O�~��D>�˄*j6,�I�go������Z�M���jjj���$9�QYc�v��o��I���5�dL�B"@Z-�C�Q%IWv�>]�[���~�B�I'Ay�oG>���;`�E��E �٘��3��׌���k�z*s�婸� $�:���j�2�\6�$L�
*!�ٰ��:�w22+�֌��O	����'���|^���̵��5a:�b�H����DD��}������JS�j��,�T��~�ߴ�\h0a�D��&i�
��:r�pix�UO5wy��@�.�|9cB~��kX�	8|�qe�w�`g,�ڜ�	��:��i]���+��Efs���������fm	��I�r���;XPX�8�,�E�?g��$��ey^5�Z���iʀgΊ�y�2͓q��$V]�����y���Nw��bw�)�+t�i� �~�egx�C�`Z:����?�j�D6FO�D>�.\v�4N9�h"�����?�7*�%��8HD��l��z*d+?{|Ԇ��i�֫��W��.�K�b�Y��q�C��*��eS��0�$�'m�ͨ�%IOnE���7�Qٻ����n�T$�&[��8��eı.��������qј�m��+����i�`0.pJ�W:M��	��Rɮ�����u���ɿ�o���z��nO�î�,����Qa�~����cG�qH�kȓ�fF��U1 �\�g׾�,�`�?�c���j��Z!y!���?,�'�E����
3��y�]E��C��	��LD�3aRK��!��];�L�cT�����F%nr���N��.E��f�kc~-r�qo�%���B���l�%@�,9~y�Sz��Q)���?��fO��ϫ��Ül5�R��������Q!�p[��a��a}��2���W��pa��g1��߉�kc��Z:���cR�qI:D��?2��l���M�����~��eH�i���F�w�����qB@�q5�ĀN¡vv��w2�:�J��"V�&6�����]}�SV�E`z��TM_��`�����w�|y���L�X+�#�X ��4}>�J�2P��M�<�t�J��es�`�y4���;��9�f�C��ӱq�F�]b��{���[����x��F���a9ly���h��;�l��(�Q_ɲό�e:ܣś_nnV��'(���z� ��6E�gTW��f��H�Д"\�m .`U�6�}!Lb��[ UA}�hQk��ܟE ��/�߾�;�T��+�C�J���F�%�n`M1�Ƅt�mK^���F��O�=r�7��V� �I�9�FW�&V�Ç3��c�&{��$Mc�gd�N4����`�8� τjO�]`��Exo����9D������a��{�2JP(G��7�RL�]{RȀ���>f<ς��#&7�J��?�G@T́l\���р2��M�9��8�٢VT9z6�	�h�\�q)M��Q��f��P��'�[ޣ$\c����I��5��l��¡�|��2����D����`X��pJ�O	�Qv��X��t8��I�u����"�^�_��x�d���X�)>|�*��M�zP�V���ƾ�h�C�)�,����S�+�ٸ'X�|�=y,�=�|��#��D��M�	�����f�/L T��G5�_Ő�F�����_����Hպ��i�Z�Q.�.�R@�SB���ᠾy@ӑ<G�����4�!����ܾ���9b4�SR���Io1�J���	<;�%���(��)X�aE���gVKJ�-T��*�9}3�8��g�����<���Ѻ����b���օ�<ʬo�aD��)���pw�H�£���b�>�������w��8WS'�^ү�l�����E>���J��/�Ř8U�W��+�9���`����7��(��.Y�L��$�Y;Z�n60����+�x��ñ�i�ƚ3�_�.��<D:���X���S�ܽ�ff�qY��e�/���0��^_+������W�?�"�:�F!GT΀�$��������h�]N�aZc�LL������\�Zc�������Z�I%�Vk�z���
V,nnn@Z\Ww���Ŝ��%Ay L��=�p����8�q)M�<������RHT�g�f 	zr���>���(���J���]��Xy��ɝ�H�#�94f�#h�W��j�#o�Nؽ�cF٥s�8u��I�*5���Y���Sx�k�%�*�ބ���{Y�kG�/,b�W�v\Hq�X�1uf����<����
wo0�z%���7Y�5E�kL%�S�,�;����-��m�%��ḳ%T��	!�L�7��um�WCV�d�dп����?I1*<u���O�c�CD���-R����� �П̑8�)�]J=;�-�O�R��Ezsf�Q�ݲ�ӵ�~�'6 ��ulS ̾�ٻ��p�(y����'f�f��i�yY���ԣ��b;|=�DF�������%�����v�E��'�m%�=���ݺ~b�6�=�O�lv�~��vQ�'���ԉ%�9���үz�a��nJ}���a*FT��9a���g��C�m�ǐ�d�\�a�A�ӏ�r�����źz�&Ů�Q�0�Six��5�������+�.�ez�m�h��ak�Leu
aP��؏���GBr�5����}��W�����S4#T���f��6�+�f\��tV�
œ9;����5�_�h*)�_���9t��<s��/��	k������Y�X{A]y�F�e�1�Z2cjz��jеchy�����=ilj����� �%��&��Jz>{�����O^ׄ_*�d[��_�J^I3�w,o-.��d�ݔ�����NBh>��^_��y���a�l|��ęx�]O�"3�ϝ�ɓ��$J4m~i_�;�$ї�B�B�N���`r��4UX���@8���PǚGMNM;;�G�h��E����k�,���z�?���y�QƖ�+C?oe������p�Ӷ�G^o`�E�4��R�X�m������/q<0
ᕀ�$���>K8rLF��e%aLĎ8�;O�[���#�j'�^�;�`�PI` D��8�$n�Ϋ��:L�Ҩ����t� ��d�S��<�z�NK/2�s���o����t�k�J��(I�? �� ���dј�Y�c�/���t�p������`�E�xiC�9ʯ�a� ��i/[��]�@���W�0�,%�]}}$jRO{�r�I�c���s���eH�d���$��yg���/XhD�*d�]8!����_ ����Hy��w)Po�tG�{)ݦc�ٖ��dֹ�뙱m�`�v��բ����=I4�Bǈ"���e���h�� +��<o����_����Dc�=pqHSE�ưc�(�˼@14Yʯ5*VY��Wl� �}NlF�9D�y8L*V(P ��w=�9�͊���b<{��UvQ>.�-�bsտ0�
l��Ҋ�;����<�g��\[ �+�t��zJ�Y�E�PO�1M2��D��͊n0��3oS���d��B
�g������nt'��k�9�Υ�Y(u���$��kv������"L�m�.9�
I��K��|�2e:�X/&z�7��L����^�������&[)���((��J3o����=E�q*�A���._��Xg�+���u��&S;�65��۷-#��r4�[gf�'�
�G��2�7\}�s��d��V�7c���a5=|y)��&�ŏ8�b�q�)�K�Ĳq��T�#������4�G����0���Qu�bt#6��ɪ��I�ؗ�XX�rU��e��Xà�1�E~�?���B���/�5m��y�]��l:F�N7�as�<����eY^�^�y{����>�	�ɍz���-:?v�]2*����M���Ԕ�ͱթ��}�j�qOyۃ���8���1{���\E�e���=a�1Zxï�-�!p���:9\l�z|��r����ۧI�@�I����(��J�]韯v ,��^*�o(T�I���V�(π�g��%�P�|������n��П����ߡ����2RJ,�^i'h�|�����)I�ӕ�58���Y�^��� �V"I"��* Ό�N�?�s��:�0F�ɳ���յ56�w���>���RtV,?����js/)&�^�s4�����*���x�,�y�sLot˦���OF���b\{@ԶL�y6��G��>6�Șp�n&���{�T�0�ؼ^��u�gT8�=Va.��o`���+���%1̠�n��F���к�̵�v},�)@��^�}�X+�����i�S���/�$���x���>G��������ֽ9��_#K>���f�j.�!y�R+�B��H_P��2m��a������� ^��T'n�>�1���	C�.��5'�p��������\�+�i��Į���n��Nv�-�s��f��W�ѥ��7���
Y�` ���&.��]̑?���@������ ;93��i�rr����v2$�^2�M���(���+�jl6a�kaj�$�Q�܃�Wg����%���-�'�P�;15�I;w"{����n�g�|�v����I�!��G�:��[ f�`�`���0k·����ku��`��ES��i��@Op�,v(pЍx�)�a9�n�:����a���Z>AE0�:�Q>+͠mϚ����B��[u�����^��r)6��b<M���u���.ڵ�O~Ȝg6/ް}O��E�#|%�k�܇�� 0�m�Kߝ�N��w�U�%$Y�jq�f�����Y�p�JA����x��ʪ�e�d��w�ٖ��4�0�ˊ\<w%/��eH�$�;
�ea��mg��-���F�_h*O��]V��63R5v�x�ϣ��M��sU� S�]��̓���%�9c�b\�_Y�5���IPp��4tF����.�{��bL�Jfy����`*N3ӱ,���n����Ӌq�v[0P���Y*�~d��[;È���2��$�f+����y����.�$�d�+���0=M�(�a.�¯�A6CW�T7O�^�G�ݽBB���"�ҨI��w�"Q(�o �f9'�8��F
���7�E+(��:�����v��:>p~�Ɍ�'����?	[��qj��C���gm�-�2��q���*�GZP'��e�B?��F^��C����vV|�z�A���sK�b��D���~�}7"nSS3ͷ�+��:�V˛�7,�S�A�}_%L�==�gN�������m��{�BS��Lg��K�G���N�u��Vg�0��kfC�h�/#S]�Y�~a��6�(ɲ���O�>^����dm �䤤���Qz���0�y�Z}��������aI����%a�fk���LP�ڣ��7��5QP��G�
Ұn��Q)�������V�:���H��3a���?$�x���A��=O������y	5v�
�tuu�i����;?�)H��:�h�4�����c���z����D,����7��s�wN��y�x}@�a��jvZ�
	���!�$"��l`m�R29V�U��V���LB������%�d+�����⣏K�{�R�RF�� |
�J�T�3)xD�\���u{�0]s�+{	��a�k�����=y�!n��Rc��rh4@	)W�*�kkO�6������zJ���ǋ���������1���v��N+��Q6!�����K��#G|d:e-���o�T��] Ч���?��ex6��1�m�� �ٚ����eS�I����֤:lKA�=�P�_2��Ѿ�
.�X#��m�����X��p��T��hŋx/���=D:�x���J.����>7�}	x!(T�ޭ�:��>�lh49��{H��m���z�0�w�Zv�:�u��a��s�?�?� �CW>�y �ˠB"0n��:F��W�EF�ɚ��C��e��d�i�~�X�}u|Qݴ�4�q97gԮ��v��LT��_L��(6�8�k
C[��!o+/��v�v=��S�'�M��t)���00�h���[���/���<��"x��TN��MtmM�k�r����$�|���C�X4:�;�-��TV)H+^?�{�~=��t%ؿN�k��P:�d��H�z�n������rH�;�c���5��wϯC۫]@�z���t�;ο���ˍh��l��<��� ψ1�_B�ª�[�e�FU�'��^��l$?��߽%��xx���'&P���H��e����W�F��+0����b� ����8��޳ֈ�Ѷ�?a���nX^i~��cM0n�ǐ�ʡ��������{#Hټ���u! م씱����־4�'�N"� c�4�����po��Nb~������WXXZ��w����; �Zw���o��r� c��,��<�j;�yte��9�?������У�|Q|}����I�ci�� �Z��F��*��V�i�.t���Ԑ���Hl���
Ǖ���S,������w�@Î}1�ay�豵��T��lK��n�����If�g�
հ��+��nPڲ[��b�+$$��b�|���d���Է��C�Ţ��2�dS�y�£y����"ً�l;��|�E��hz�#���r����B&5v���kF�-����*���*��dj7!����L�]��߾���'�9&���T�xs!�l�3%!��9�
e�tPE�7ʂ���5s�\ل?z��1_)�̓@�����34��E�F�M@F�V'���^#�����I+�.���,���(K�x�$�&+�w1==Rhf@\Jg���k5,�)**r�/���%�O�]"�C�|�M�`�{���(��+�#�Df��W��룯>�g9�^���SƲ������k5��75E#�r]P��o�Mw-��W����Z��Ff�E�6Jx�Ei>��U��[�ˆ�!I�O�`L��)�^��or���R��11���6�M!7h+���㇍�����!��~�7�{�a�o�T������㖲|ȱ^���{l�=��{p�	?	2�.)����r����%s�`O3����̒�%/��~\�l��y�����Mvlc��n����Ӣ�"�ơ\���c,l@�R������"2H��|��E�&]!�� ��x���&�g73�W]Ᏺh	�~�K��WzF��u�jb�+�)��.]��w��g!�X�#7b�A[���'��w�����VT�2uɖk��c���eq ���.*Y�:�0��O�1Fd���ݾ��)<�L��%�/Y�.{C���(�4��$����F���g��P؝P	H���6@�J�d��6,>��~	1��t���́�j U��i�ʅ�6���U���i�e�Ŵ�	3���4��=��!N�O�&AzwS�6g��B�2aW���eZ�β�ie�O�nz,mE���#�Y��ݳ6*�e��~��[�8\6�! ����#���_���O���T}���g�����y�A�����z�.�v����/_��S�B=٭����{ IH��m����x����}^�CQ�h�?��M��h�r����[��=KP~��A�gT�zxzn��<5$|w��"��|���lV���吀� tm�.��A�4I�ݫ:7�fۙ�K[�ۯ
�/p�O�|#���2\��|�b8t4���Ό�8���+�߱��V���e���T���F1$��O�|���P���+���ݐ~M諂����qI�D��!��O���?od����'�:�\E�:�~(��*����v�<a����v�f�Z�"GEa�5��v���)��}����:!��7f8	����&r�Ҡ*%^@���z���Y��F�s��(��Zk�IH�㆚��˰�J�����tR��(�ǭ�T�ټǞ�K���ǫG��R9�����[�_ʯ �Pw���J*w�_?�~�Ɯd�s?�gS��Z�|�^�,��`�����V34�p�nբ��WB{���I�.�����l>Z}�p3V��+�w�<�5/�V �~�]����m���{*M�WVS��3�ِ�Q�)��#E��D�q���E�i��
�:�����Y��lB��^&�g�6�p񐑌�O�?h{-�'�<������qZ���f�uHqS�9b.<���E���k��;�A�G5+���v�Uí9>�$�,���g��w�j(C�g4g�j�7�֑*��m4�%��o���Co��"N~yE]f	�~.��xzO5�5�k�G��Fx�f��V�'l`�G�5f�V��8��?�.��3w�@2�Qyʴn��M��Q��/z��5�I*jwg����C+�
��-�#\���X;�$�8G��cb`���T<���Ҭ�xL�އ�h菀�̈'������	�;�;�y��i*L|SLn�;�	�v�٢���0�M���r@DA�j
֊c��uy����j�Wט���
Sp�2 h����Ꙕ�
����c>�W��I!�\Ѩ=���FB�y���*P3Ǵ����oiS�2��\a�Զ�auk��)�DL+�S^|N��3�}�m�"P�A�D�n��U�3��cx2_��g+(�[� �l��h��jE}�G����V&����R��q[�����L����ڲN�K���K�����c?F�oH>wRM�t�-�-
�*�nL��\�v�Ki���dgX���cW]�]�,_�Z+?�C� �F��7��=�ou6��J�3�ćA��HC� ��R0��x��#�l�S]qנ�Jߞ�)�+����ھ4���d`�xmO=[�������j���}��4�(���b�Y�t~]�f�ݧ��cLp���4�Ϛ�P�ElN)n�M��8�'�%�-O�Ɍl�1�2w�uk�����P����F��_��
��KCu�C�n�Xu��1�'v-])�ޗ��H8$�}#��Lm�m�#W'拉���I"[R����Tx�>��K[�÷�Ȁ���w����$4 ^�rK�q�
�g7���2�.�xsa�V}ɼry	�"�qg��=�F�Eߺ���?�������YD��r�Yj��EO���O�r����[LR�x���ș� n�/Y���Hro�C�y��"W(N�N��YU������|j�Ё-שN�U��fl4�qlb���R�ԥ��������U�4�������w ֎�K�����:v�SG�`������y�`-0h�.`�b�_�K9ߗ��pFН��R�s����X�ȡ���.�C�=� ��`g� e���Dt�l9Ll����QQIɫ
�$�:Tۚ��u�C�@�D��sD���b��Pv�=4���y΁�?X@�"gX�*���B��;T�m�(0reVn�v+@搹��%$<�k�=z�g������X�a,ku��?�k_mLi�hI�o@i���Q������ņ;��0
B^_|��H�K��!�+�e��e86�O\c���B�)�n�N�#��!����~�����/0��D4����:�n����@K�t�.�Yp_��ș4y�B�$��J-��������>s��y��SNßE�En��,�r��|5����q��"���&'_���s���f�"�yg��y	V�+g ��<��D\3�҆�{"��-k�����ӛ��HGs�Y����A#�t���b��[�+����mYT��j�b��&_{��W68C{��u��%$]-��!9�,x���A�E�F�{����u>�ǉ�b�	���������_�-c��U��x.`vP�m�򖚠�qj>�}mP�d��Iw�������ٳ�6���X�|4���b�o��8���ϥ
h�ݷ�����d�R�DQQ��[��C��h���d��"�ӆ�lU�?�~%Q��2�W�Mdn�tz�f?��F��2{��b��m!U�J�Q�3Nd<��Sb7�:���lTӦV�w��n����1���a�����k�į�5p����< .�w.���d\�L��7g����Y�6��X{�P����ҹ�uo��;Ȅ�|]�'}{��Xw��R��d�Kۢ���P�;S��G��ymt�F������#�`�b]��Z}��ZU��3Qv�&]�Jk'��cE���EQ˴�^�.��>�F֕�ʙ�Q�o�ɾ�R��>�l�[�kmt�.&U
z[��M"��biJ:f��~�9�k�O���R��
�ܘ0Z���3�Q��3]"�Cr9�*0�*�/ʠl�?{��*F*��M�P!u��,S��ɘ�Ed�I6J�����{��=�I�
(!�-�C<?�w��Ut���Y������UL�y*a�9P�����������D�ϗ5�a�T�O�� u[�{J1�F��' ��>��H޺�ƸJAA���wv�ï��1��u��/�$��Mk�A!KM�*�Պ>;��aw��n�Q1P���%�3Ɛj�����ye�G�6��}C���UV� u)�ao<$��������U08��c�
���N����k���xk��0��RSv�_��{���W��(.*$�WVbT�yx̍!	�)�0�t��84��4�i����_�fN����=*#��مh��ݯ\L����2�W^��_�_��]��̽������칊)s)�ê��y�C�����D�V�sR,.��!��ۺ{d�<DK�2$��&�UM��<�\{������Gr%��{�ٵ^\��J���h�<7^&�G��H��o�tm�SQY��k���G$��M�3��������]�k5��9�~t+���$�hU�����x\����Q\��ЊU��Z�JO��M��禡�;�7��j����&�4��(�j�u�`0�Q�j7Y�t��t��]�A?��7A��Y�Wom<)p���-ԉ1ެg.�`#���S���J�0�c��C"L�֌8�bc\0g�2C@�a��%��^V��.I����ĕ0E2��n��[��C�w�D�*(5I�f�(�S�"n��iȚ3讠nUw�[�;7
#R$�}C���b�8,��E)}��y�!�I�աȆ�J��1׌e���biׯʤ�H���O)4�j�w�X�qxʧ����g�-1���ԾKu���B�+�4w����������t����}�̡>�<�P�)�)K���[��	hb�G�"�D=��H��M�y���@w(�$Q�Z��K&�-�7Ny�8FZŘ#���R�8����9b3@�
%���F7�
\��Ch�s�eO�0`���i�e�����ϥBx���	�E(J�6�P���D�3d��HPI�j���\��F�I�����m,��L��1dwIn��w
�B�d{I��=����2}x�:����Xjx�	���f�j�/R5��������kjbC�F�:
�.� �ś���A3
�����"�-��}&�=�,#�'��k*V����1�
�@�#]�ab�Z>E�
<c��]������5)�\`�س*n��Gm�j����<ʽ
�9}��&�l�`����;0�*M���n�'xz0�Eh�~�wS��I����3��������T(m�#��9�j,�O��jN�w��I���
��|99��d]EĿ�r�o�dT�9�����4���-U��l�M!��&�ґl��'��*��)8��2���͓a��|�&�n��ڼ�dP�_�wB��������O�>���W���tO)��"S��+�t�,��K�꧶�p��R��	%@�ww+��bŭ�/)N(���G)���V���=�_63;��w�GΜ}V��F%]�`u���!�k�^�i�Pnf{_���9��]R,"8�u	�ʰ�`F�Q;GvDً���x��I!�=��W���_�6x,r���mBO��;]��$��`*I4�����_���{3.�"��R~�L�O��fA��큄�~���A$�$�,ӇeK��[W����:���g�8l��Q�L�r�߁�~wL]l��Qi�I���,�^"s�,�F�mgOY͸5�~x�6+�ڳ�f�hă�>p�H�@��¢i����+q%rǌv�$���Ɖ
�W�9����n�A5��)��?��M��� �}w��H�;@� aTM�< �]�%fS��e"��6�)��\02�:e9��?�jEP>�o/j82�M�B�Mfz�:	��d����J����ĸ��9�sx�-�|��\�75(O���c��@U ��$s�T������V�O��\C���U+���V.�c߶��-N�I⛓�V���7UMvE���e8��v�r�wSR��_�P���yT/O�d/�^*��n5І�4����1�u9~���'�4��ۚ��|�4�m��5_W(���f��}�e�ok������|�x{b��z��E�ԱZ�z������[mX>Q�^�����wv���֓V��$�_f���s<F����x�vH5ZN�9���g�Z�XE��G7���a(��_�B�6hF�/�L��8&�lm����uWβ/uME`�e�$�����U@��zՂ,������U3
��Ɔbjm��ܰ�D�>��*ӏ�&e��m�W�T$Y�W��3�]�DZ�V]$�� kQ����[.cF��x�\��Re$��2������
�R�k	�����#'M�a3-��?a�m��?�HYrA�a�g�S�c����5N	5I1�td�ZR�AX0eh�<L�#�a�g��p�pgq��N����ف�ܭ���g���k���1�^u��4�-�\~������Gf]���$FF�����́�ǩs��y�Iی�w���L	����g�{�Qt�֥4�`wty
+��e�sCT]�Зݦ��+��v�A?���nSXpJl��`��S?�8@�sI�>�zK891t�5��m^�������'���22�}���o��:p�Q['��^Ɲ~)wk#�V�L-�?�po���,ݟ���WQ�'���j�U�A�4y�<oq�҅`@c��1���8��N��-�#)M:,R��]���)4=<�;���ا�H�՝�Fo�Nt�+Jv�����c���	�vO�����Ie;�p�f+!:�����[�̫ �VY==�*ӮS����@QŦ/a4Z8c����l�Z�ʠn���Qm�D	��/C�C��-<�iU����h���Y[2��H�U4���wv��Y ����,�җ��/p��nɇ��<�&v��i�"�3m��d����,�Ȭ�Ը�3[���{�mUd�*09R�Aݔ�GI�P����.�������-��?�O =�=�}��f U�}�r�N�|����T�D]�D��݃.B##/~6�;.ߝ��Dd����z��}�A�M�F�0�1mr�w��`쿪����0�u���I���:O_tI멊"�}f�w�t�"w�2h˯"���S~�v�m����>��#�ufK���=���Uf���ǟ�1�es�t�Q�)�����W	2��w�)�� `؇X��ɳۋ%�w�5NW
2���vӠ�f^�^o��(-��+�jܳ��|����"�I�����qBru���>@�X�P��4�c�(�L�V��]/�p�����x�8M}ٗ���t������D=�R�SO�Q�M��D\j�Fm�cɻs�,�����$����H(�̱Q�}�>J/#g���2�
���:����������(v}��ҳW�DU�Q6�&�WW����!{��A2��r0��}��Ew�5��o2O|�R�-���o�t��1���@/�]�fӬ^�.��L��A!�i����X����P!I��Z�d$4a�gd%�W���O���=z��nt����m�x����-т��ã�kE��3utݤɥ�-���>�҆�0�;Y���#B�02%Kڸ�׼�?<
*۸�@Ϻ;n������}����uy���my��ψ3�v�q�d�Ӥ�[�s�4����_{������lN~j¾O�]�u���g �$��C3��2�V���~��1φc����L�)ޣ���`��X-1mF��W42�8	z|��'�N��>@�k��+�:Du�/����k�Έ:�z�Z�oٱd�l��Ǵ58Լ6z"��ì�K�t�ц:�+��Y��v^b9~d�߼�{�?�7Q G1�M�5������!�L�ļH����N�P�ڼֲ`��֮%��s�ph���ҋ�>�C��Z��������y��$5DOGZ��O���Q֯�X�`bF0�o׏�ȓb7���>,���ٰ���#���!�ss�Z�o�1ӭ�Wt|k���{G�����A��H��j�u�0���8#�*)
l3�'��
��[vk1ۑ���n�|��tH�N�8�|��{�٭��eFՃ�x�O~���۸=us�D��>�_%�(�*/V��
fPҷ�*��"W={2}��Sܵ��v�YWt<բLq��v.�M5�������t{wT���͵Mp��S($	į$#Du�w�v7��ܬ�v��fn�oAw�H�=A"PF"f�a�����k�gL�h�DX�l�
��?��A�$�6]� ʱ�AG& 52�5Ӑ�,j�0.|���y������R"V�quGe���xK
��Q�#6sF��`�ܐ��X	 �I����5*_ב0	MIF�=�X�]c�"6'��G[[���b$�_�#?"7��U����:���B�H�������e��d=#�>ܞV�W�j��D�Լ� ��	hi��k�)�Mż��4!ݭ������)�rţf�2�h�&+4G���k�8���v�<��f�@$��>ו���=O��u�)�\��[?�64���P��iQ��ݲM�I��<x#��{o%ܣ���[&-��i�rY �� E�X;%嚋�t���?J�h���B9���TPR%R����{ĲH88�ks�����܃@�f�0������c!�\���-����h*d����M�f�ʾ��kThC$�~��uhD��~�ܻ3=�4�<�� �ANW���%���~aN��DlZ(�rI�B2?�f�ߋ�]]�8�`���O��w�,At&�>qR��q �<�cJur�-ٱ�	w�
�\�}`͂��-��蛷���+>.�D�B�1eVx2���6�vY�2N.�\���r#�[]]c�2���B$����v��yT���wXA%���,J�.B4��M���t�ш�@~Z��3���.�v�qx����_����D�°�YY�pHR�}��ѵz$��=�p�pF��œۘm�����k�D$�K"����g��K'p��/	��G�?���O�LW�Ѓ��%� 
���v�	�V� �\�\�[$�0��Ƃg/d�����ˬ�5��=��Pģg["*>�ԌD��Gq�	uou�r�qV�lQ�߬8֥�����qrJN��ۃ�T�Х��aX������)��[�����Œ����H�S��B�9�E���5uڈ, ���DZG�8��.*�[�D��_�X�+�z����3k$�T�O�����Œޥ�y��{1�_^�X��-ZVƻ5�s�}#��!_&��'�����&;P7D)��玝?�9wvv�(\�v%�\?۾y0����*"�N����V���q������-$�`/xC�� ����W�M���Y9������_\��555�
��2�}w��ǰ4�D�=���U�#5P���'���K��V�xR�ޛS}��!kd�V���&����{�(�+�΂[��E�]-E�(��ռ�Š�!H�W�4���,�䭵f���'-Z�PpK���%�vB�=���^�|�/�!!�HG;�G�``�*�����+[R�7�	]�σ�	�:0����|m\�(H��`XV|;?����a����?x�0�K�����}Iw��`<G�lq���A��Y�8��l��:��'�r���1E�0%��DMvfꘝ�H�J*ǯ_E!�@��|q#�3���8u9 �]x>њt�O�׋"�G���GeD��B��5��ԯr3c�\p;�� ~�vF�Ɏ���ԶF7+�~mĨ���=Qɻ>"I�����e�����z5�#�6�ip�G�@5d�u�z({����2N�<�ٔT0A��2#�K;�W��x?����Fl���cN������Wn��+�s9��I?"��?�D�k�r���{��*L���뿉�Ī�av�E�{;T�$��):��A�im�Ͱ����H��w�uK��!�c��9娹d}�����O� +r֛r��o2�����;|o��Z���Z��XLV�=��-����1�ׁb����B���ʿ_K����\��S���Q��/GM����˄s�A?%�9T��ȹړ���Foļ=�6-bV��ۡ����
D��&.9T>����S��N��Gl��Z"���He��2rz�4N^�wN�
��D��r�9�E����ߔTTT��d�%w��Æhj��i���S�j*�}�+���L��%�g|��xa�'/��nvR���O�@y��ң1����+~骥��k��ֶ�b	:$@]�%��Jtr������5G���FǶZ�_���3ƜJ��Ͱ\�[�@"<��3"u��)l��+�v�U<���?�qZ�/Nr���{�be��b��%+����0���S4�b�«F;��HcE�k!նs�R���%��X�-
�r��H�oW��R<�b�Kov|u�eK�+��̃��ZS�nűy���c����a��Z�Ϝ���������O���رu����X�2N#}L�6G�쳭��'	��0�� 
[���J�]8�� %��U��7́�9�S~�PF7io��<dPۓ�6�%���n4?s� 暭a���T�'-HC��[q7bQ�T��g@��v�Q��U�P�dH�e�c�����j:�%���渊�(b���>�#�Bë��Vev�4�j�A��$����j7!���gc��>��Ϸ��Ѩ�B�����U�?_��#Q�PO�{�ʢ����K.��gʑ�4"u72���tL%�����t� eH�+;ZCj��}f��kzE� D�TT�#%r�����tU4bҊ�P�D�V��+�	�+�<�"^�s��H�Ƥ�rֻ�۳�VaDw�q5���(h�k��n݁W�Z}kW����������/���]$~��nA����x����޾������ Z7a�t ��Ո�-~�0�3�o"���)d���)�.��[	{w��������bL�J�A{m��#N��lY����4m��^��M���LG�J�>C��|���2� \��S_�Liey��ј���)�
��;pd�A��U+Ig��q8���Q�<Րw��PS�y킇8����D?hL"�4�k��d�2���u>��R�+��Z���#�����c<�A7��U�Z�s�|e�_�� g����_w�*ꨌb}�!}�z��I��ϧ�mȿ��\&�a!�iY��".2�Sc{31TN�E��6��Y�V<^M�H3��cߏV���T*!�"��.�֩�F��������QVMB��^u��#ysŬ���@��z5�V�_��ex�f8���t�WXh~5xG}��N�CKl+ 6��C?
���!��DmO4W;Ek~�/�����К�"̨����杁��D���=�q	�,���v��.��"��N����葔�ݻ�3��_�F �������AFV+
��w��O�ۆd�R�h�F�5Ԇe�h��yi:�8�	Z,�xQZ��6���啧�?ŉv��"�4ٷ��J�-�32��N�}��0����l�/V �_r�|-���,���4���H���D#�)��R.�Mn�>?k����/��G�Q�*w��R��M�M�
̖���#��q1?7�G3���Vx�7�aYt� �-�6o.�C	r����ΣG2
�rO�x2O��]�?Oo�A%�f�t���}sC�=:�FŔ�|�KYg����YV�pFգ���yA-��+[}ѭ&���?o���5�oi:Pch���.+䎌��k��p�A&���*gd��O�H�f�>��x�q�#�@0�=����]�¥gХ�*;Xۜ7��j�)s�5i�9j�WvY���tdt�_1Xno"@3p�\<��'S3c{�5/o�j�����Mj�Ol����<8��g�<��{��t����/h�]����r��Y:��A�q7!w���(�	z�Se:1X5�-�O�^�F3`�r}2N��o?\j>���jl5NtK��������z<�:��'�]�C.yh�md��0[��WQc��ZW�rZ� |*�g��*e:'�vɰ=h��#
�͊{x^ ���*Q��C�m��p�����ϧ2n�m'ďG�a�M|��tz������,;�KnY[l����\©K�t.����/���!a�Fbت��O�\�wE4o�څ�wiUEl&�L,%��o�8p������kE�p�5^��L<�G2�Q{-�����M��!�j��Q�k@-層d��ߋ��U%==�F�GsZv��{�(K+����t����h�-����kAu��fe$)�.��='9��!�%���E�݋�#�'���%{�����ߏYā��,���uK.�@t�C�|� ]�(�.\ǣ�?(v�#��/!7�&S?Z�e�9���]��?����.-4����/�!7/�������\��	�n(K�X	�e��ku~�@����J+v5�ǭ�	~z��Gt�:U����Z��u$9FE0�}L(Q	op��U�)� 	ױ�0�]�'T���h?�o��8K!���^w姟r~������������V!͐�k��d��쪸p��#A�/VHvh�*� �)���O��' ZB��HWx��J8���u#�%6*��@j&.?���A�}Q�0�����5p���i�a�Qڃ>
B�G�����{Rie:�l�������-ى�p�aHT:ˏתd�đ����է��?-��Y[�m�v�5��K�� p��<ҩ§�Fʾ�y�����zQ�v�8�&ii:~��
�ri����k��E���p�fv�r��lR[��?��H*�R�� ��þp�y[ә�`%���~�lNu�Ge�O�5Z���%o��e$����Um���W��g�7�q��gBY��^�QU��)�]���|�K�)��H��t�ع�2���o���r��`��}ZJ��]�	|~\/�~D0h'	ae������sjfڎ���D����u)�?� M�r��a��\��������9e��z�3L#AAͬR�x�!�T?LmЖ] a79P�e�py�o/ڬ�-|�ȡ��4�5:5+�J.�2�k4��)Q�����,��㦿�i���9��}��VK�B����~3 �\t^7�]`��@������,�2��.5�$wa�����[�����#��1�.�d���1d�"��0���~xH�w��i-P }o�t&Ţ��ߟ$�n����e�l��z�/����z�}����W�)��?a�s�/s���D�hQ�L�J$���VC+".Đ_U��}D]g��{�1:8$T��� ��Y��*��H�8���>��������	�=o(��K�^��٭��*	��m�ׂ|i����,Z�K�͋��`��DN����'>&�5u�n%�{:V�fa�&B��b�L���oT�]��sKHhg������^�5U�I���Xa���������G�h��t'����Ĩ�S17?~N����fq�R�\���:-�C����Ո���J�5{a�E�X��@�a�2�+�0�
�����t����
p�9ɻ�3j �e�{��M�O���Epr'1���Ma(�L�x���b���Q:��x�I�`���գ)Yv���#�*���ѓ�-��^}
с>�R�ˑ׭52���k�77�'���/��C�bGj|��F���8��sq���d�����z�^q�_l�?v�FZzƱ�|��
�ھXG�Yz�1�|7C?p��7�!��&!���(�ـ[��B�.<��'I@
���3Kl.����e���nG\wd4N.��#|��C�`��z������qæ�W��i{��bA�T��n��d2�̾�#T��ǴwAٰZD�xG���(;����P��)]�,}�j��Z����NK�Er1]t9b�����!�DOO�k<YTŐ$��Y�#G�ra,jL��zF!�.T�E%BV�g%�m����Vx�,9�X~]�G�G��QӛJ������;0~a�g�T�ѵ��Z���)C�3��d1�N�h���k�E���F�(�^�������c�␮i9���WO��&1�ڙ�e#@�ű���������+i���WL�H�J�<�!S�o<,1z�8ʋ_��tఐ�r
�1��X��(;ͫ�Cz [�>�c��HԸ���eU��N��lF9_��Z�k;zh���1g
��(J���l�p������m�3����{;�3
�i����>3�)_�m���]q�<��ح�MTH���r�.�oڻ�j^L��&������#X�)�9�N��Q�k�"k6�ܸ�3�i�$��e%)��n~�� H+G�3%����� � ��A��R+06ۄ�i!��j:�p�Z��{�.��NRuBVS���>�׮��5�)��ާ�e�?{~|6y��ꚫ�7�F��פ��hv{�&Yuxx��Q��^��jk�4����m�&S:���Kj=W6N��(�l��� ~�KX;�ւ�2��#R6S�M8M���Pm5|!��^
%]�٤�5y��7P��-���g{�������4X�*��V�afG�CLm(��}���k�d��F] �5�'�s�'�	��r��]�,�b�k�8��x��`��ɿqUFu��vD4��/��=g��gO	)�x�F��T��p��v�2ʪ��zע�->!�25��k��ԁ�B���
�T�%@�'[\�x��PM�����3�v�x,�q��R�zK#���I�^@���TS
6�M&�J��jF)TY
롧���0�k��|�`�n}�a���	��ۋ4����Y�����69�
��,��V��"�9en���>�Kńde�>�DQ4'O���9S[���'F�i�A���^�~+�d��S�FT1�<G,���xQ�f�,�N�Bs:�]���bL�"��ZŘ�ƊU�#�h B�:4w`5:В$�,����'t}�)ԞF�&y���aІi�g#h������_Y H\XӪ�|u{I�H������kh� �^�X:�xg�e�1�տt�bR���
H��)�\�elD-��$D3���(�|�N���[0��f�-LSg��P�}���+�[W&g՜_G��訽�X`�RL�e�SK/C�gf�~�ư�b�6����u*48dU`�}j��~ؾi~5�:� ��7ۛ���	��")=
�F�p�&���<�|��+x�k��B|�
�u!W�l�o�u�}�/�j!���٤I��nԴ��=p��w���v<��N>/�7R�~z¡B[�3�z&t/��y$�A��������{$yB��&�����������D�����du4�ր����pZ\0�^Ct��
�2EN�
�o>�E%�����r����p?6= ����sL��ۙW���smu�9�4YԒ���[x�|��o�Bo�����?����iЃo)y��,�	x�td�𑖍��8.#���f������V\E:�J��������d�XC�R�N���\Z��͕��#�E�m�M�#�ō.y%�#e�z�Xa'ߢ�~e��
�����RFC_�:���|�mkd�1C�Q���33��{Az�C��D�%aV�.s����j�z՝����$�z���1�+��T��#0�r�qjq>�����f��6&�������zIR��IЋoM��o׵�.��Lcb�������i�M�W�Dv[����3��(�7���3�F%ܖ��̷�S��z�F�\(���)�!X/�8�.��	��tP�k�$�Q%���cb؇ổ���59��1|[���=�����x�gK�t��r3���C�x�����������3�ƾ,s,�5"%e��LOW�����Qq�bB�;�A����ׂ+�כ����F�/�⻍����o��P��&`��q��;`���Xp
mڌo�l�v/�уN�m/�5����؛9� �Y�N��9w��Md�`<?���� H*�����;#�����ϋx���]P�ҝZ�&&SYj�����*�caA�:�X&
K"�.i���Nb="����Й��e���n�)ʯ{g�ǯZ÷��O�/g&�Ir���{%�]����2�3����@`e����ֱ�Y|��'X�
��W��_��{��?pm\��F����y�v�o",�q�y���`��[�D�c���x\�D�Vqeo4:�l��֤h#V�f|����jy��N��=�Vl��w2U%|9a������}�[X?G�u��o�I�r�)\�"A�~�A��VϿO.B&rc��t1OX�ɫ���b"Jd��}��8.����=��5X��e��-t��嚓R��R���.*T�F�w�5��x�"�z���K>�r-I>m���I�2�̥	����BN��[�K���?�^����]S��]���~ԙ��s*�k[�U;�aX�5=�eJ�M�+�; ��oz�扭��Ō�Y���z�t�e���I��͸wt��&W��s�iQ�@hٞ�TZ@��כC�VC��2$�Ԯ؄�X�߷V�ke쥸���8����A�@���N�'

���>��
J>֎7��]FT��N�����8Dv+�"���7N"�?B�^��f���La�����Ǡ��ʂ��^�,"��"#!I$�N��0Y�~�L /%9u�i���PK   D�LU�|e��  �(     jsons/user_defined.json��mO�:ǿ��W 5������Bե�j�҄��<�h%��v!���2X��1����>����s�'k��M�3�K���$��$�֏��eE�߀tewXW�Yg_�^��
�g=�'���|f��~���,\�PE���>q��&��,�F�p�� �c�Q�e�{��0�)��Э���^=ۗ��m>�d��v�2�?�\d����6�ʟ�f�4O������l�݄��b���P�����x�ޤ��c���!Ͼ��i��+�|.��]VMu�m�a� :�0���y�����0�?��&\'�#Kd=��#q|�1~nv5�E3 +�5�f QF����4\e�&a�T�.��)#������T���!���a���2��G�BS+�h�� ��u�;��Rƺ\�یP�Yq9�nF�Ռ4��f�Zκ��(h��l�!nƊ�$J�2�_��it�B�P��=�=
��fu�nzP�PQ�w'�����:��$�E��/S,*�N�!OcQ��e�!QcQ��z��X�u=�>R5EWG|<�b�8���� Qk��ɚ�%��dM�r�#Y�i����Z�=$k��t�d}{��_J㇬�e�3�,�I�ώEpU�FEޱά&�w�w�uR��`�2'q�-��p�O[*hIU|,�#BSB�᳡1��ALl!��̇��Y���X4q�a,-�1v�F4��C|
!�^�k��~&?H��E�u���g1�c�J�,܀I����O;�T#(	��BǛ"��B��Q���o�P�&�܍b@>�e[p���Mb��8Y-� 5����36��
qhi�CHjq�Bn�U%�Ʊ�>A0���/��7GV��8���PR���1"�♺)��M�CUpI*xC� ��/��ٛ1��-%����[�o����.'��3Ū���]�?:_8��K �ѭ+)�	61�n=�:w	��eE2�4�k�	�-r���#E���.H�˞��.q�����F�{0� q��$���S���B<�p z��:�EI���n����V[����ٵ��c��<+i�����ٜ�$M
db:�$iS S�i��Kz��Wp�RҮ��>d�
̌ܣ�̵fTI;��T�)Pp�i����)*B�a�:8�w=o�h�Ao��58C��6=��Nc��X�K��~��?~��ñ���{6��l�]���|��o����vy>.�o3��H7�.����2�~8���>�V�	�4���2)��5�z���k��H��6o�� �`8��-�c;-^�4��Ц.�m7L����o�5ek�)b�i6������ʞ\�����A�0�{�-p}���@�O�����V�E�$�A3@yY����xǨ���^$�΁T��ju�7k����N>XI9
�o:`,84�7�]P�q��1��O<?�1��t���2CǇ̓j�"��.k�2�~�B�R7��������Q���j�JId��xD%w#��	������_PK
   D�LU����R  �>                  cirkitFile.jsonPK
   ��KU_�6�3� �� /             �R  images/062f1f9c-d785-4821-8269-cd0e0f0d9a41.pngPK
   �KUM��M, W/ /             FK images/88f9db7d-1b4f-4095-8375-25787367c0d5.pngPK
   ��KU�р0G3 �	 /             �w images/c35f35e6-9335-45d8-b9d3-3c107d870976.pngPK
   u�KU�b��� L� /             t� images/db75ecfa-5437-4ae2-b047-1b58b40ff187.pngPK
   D�LU�|e��  �(               �5 jsons/user_defined.jsonPK      �  �;   